-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    read_write_bar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(9 downto 0);
    write_data : in  std_logic_vector(31 downto 0);
    read_data : out  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMem;
architecture accessMem_arch of accessMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 43)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal read_write_bar_buffer :  std_logic_vector(0 downto 0);
  signal read_write_bar_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(9 downto 0);
  signal addr_update_enable: Boolean;
  signal write_data_buffer :  std_logic_vector(31 downto 0);
  signal write_data_update_enable: Boolean;
  -- output port buffer signals
  signal read_data_buffer :  std_logic_vector(31 downto 0);
  signal read_data_update_enable: Boolean;
  signal accessMem_CP_0_start: Boolean;
  signal accessMem_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_136_load_0_req_0 : boolean;
  signal array_obj_ref_136_load_0_ack_0 : boolean;
  signal array_obj_ref_136_load_0_req_1 : boolean;
  signal array_obj_ref_136_load_0_ack_1 : boolean;
  signal array_obj_ref_140_store_0_req_0 : boolean;
  signal array_obj_ref_140_store_0_ack_0 : boolean;
  signal array_obj_ref_140_store_0_req_1 : boolean;
  signal array_obj_ref_140_store_0_ack_1 : boolean;
  signal W_read_write_bar_144_delayed_4_0_143_inst_req_0 : boolean;
  signal W_read_write_bar_144_delayed_4_0_143_inst_ack_0 : boolean;
  signal W_read_write_bar_144_delayed_4_0_143_inst_req_1 : boolean;
  signal W_read_write_bar_144_delayed_4_0_143_inst_ack_1 : boolean;
  signal MUX_150_inst_req_0 : boolean;
  signal MUX_150_inst_ack_0 : boolean;
  signal MUX_150_inst_req_1 : boolean;
  signal MUX_150_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMem_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 43) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= read_write_bar;
  read_write_bar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(10 downto 1) <= addr;
  addr_buffer <= in_buffer_data_out(10 downto 1);
  in_buffer_data_in(42 downto 11) <= write_data;
  write_data_buffer <= in_buffer_data_out(42 downto 11);
  in_buffer_data_in(tag_length + 42 downto 43) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 42 downto 43);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 1,4 => 7);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 7);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= read_write_bar_update_enable & addr_update_enable & write_data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMem_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= read_data_buffer;
  read_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  read_data_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 28) := "read_data_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_data_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_data_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_CP_0_start,"accessMem cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_CP_0_symbol, "accessMem cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMem_CP_0: Block -- control-path 
    signal accessMem_CP_0_elements: BooleanArray(28 downto 0);
    -- 
  begin -- 
    accessMem_CP_0_elements(0) <= accessMem_CP_0_start;
    accessMem_CP_0_symbol <= accessMem_CP_0_elements(28);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group accessMem_CP_0_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	10 
    -- CP-element group 1:  members (53) 
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_computed_0
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_offset_calculated
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_resized_0
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_computed_0
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_word_addrgen/root_register_ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_offset_calculated
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_resized_0
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(1) <= accessMem_CP_0_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	24 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_137_to_assign_stmt_151/read_write_bar_update_enable
      -- CP-element group 2: 	 assign_stmt_137_to_assign_stmt_151/read_write_bar_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(16) & accessMem_CP_0_elements(12) & accessMem_CP_0_elements(8);
      gj_accessMem_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	8 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	25 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_137_to_assign_stmt_151/addr_update_enable
      -- CP-element group 3: 	 assign_stmt_137_to_assign_stmt_151/addr_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(12) & accessMem_CP_0_elements(8);
      gj_accessMem_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	12 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	26 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_137_to_assign_stmt_151/write_data_update_enable
      -- CP-element group 4: 	 assign_stmt_137_to_assign_stmt_151/write_data_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	27 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_137_to_assign_stmt_151/read_data_update_enable
      -- CP-element group 5: 	 assign_stmt_137_to_assign_stmt_151/read_data_update_enable_in
      -- 
    -- logger for CP element group accessMem_CP_0_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(5) <= accessMem_CP_0_elements(27);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	12 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_sample_start_
      -- CP-element group 6: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/word_access_start/$entry
      -- CP-element group 6: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_136_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_59_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_59_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(6), ack => array_obj_ref_136_load_0_req_0); -- 
    accessMem_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(12) & accessMem_CP_0_elements(8);
      gj_accessMem_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	9 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_update_start_
      -- CP-element group 7: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/$entry
      -- CP-element group 7: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/word_access_complete/$entry
      -- CP-element group 7: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/word_access_complete/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_136_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_70_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_70_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(7), ack => array_obj_ref_136_load_0_req_1); -- 
    accessMem_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(20) & accessMem_CP_0_elements(9);
      gj_accessMem_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_sample_completed_
      -- CP-element group 8: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/word_access_start/$exit
      -- CP-element group 8: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_136_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_60_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_136_load_0_ack_0, ack => accessMem_CP_0_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	18 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_update_completed_
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/$exit
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/word_access_complete/$exit
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/array_obj_ref_136_Merge/$entry
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/array_obj_ref_136_Merge/$exit
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/array_obj_ref_136_Merge/merge_req
      -- CP-element group 9: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_Update/array_obj_ref_136_Merge/merge_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_136_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_71_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_136_load_0_ack_1, ack => accessMem_CP_0_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: 	22 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_sample_start_
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/array_obj_ref_140_Split/$entry
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/array_obj_ref_140_Split/$exit
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/array_obj_ref_140_Split/split_req
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/array_obj_ref_140_Split/split_ack
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/word_access_start/$entry
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_140_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(10), ack => array_obj_ref_140_store_0_req_0); -- 
    accessMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(22) & accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_update_start_
      -- CP-element group 11: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/$entry
      -- CP-element group 11: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/word_access_complete/$entry
      -- CP-element group 11: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_140_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(11), ack => array_obj_ref_140_store_0_req_1); -- 
    accessMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(13);
      gj_accessMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	23 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	3 
    -- CP-element group 12: 	4 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	6 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_sample_completed_
      -- CP-element group 12: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/word_access_start/$exit
      -- CP-element group 12: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Sample/word_access_start/word_0/ra
      -- CP-element group 12: 	 assign_stmt_137_to_assign_stmt_151/ring_reenable_memory_space_0
      -- 
    -- logger for CP element group accessMem_CP_0_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_140_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_140_store_0_ack_0, ack => accessMem_CP_0_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	23 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_update_completed_
      -- CP-element group 13: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/$exit
      -- CP-element group 13: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/word_access_complete/$exit
      -- CP-element group 13: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_140_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group accessMem_CP_0_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_140_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_140_store_0_ack_1, ack => accessMem_CP_0_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_sample_start_
      -- CP-element group 14: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_144_delayed_4_0_143_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(14), ack => W_read_write_bar_144_delayed_4_0_143_inst_req_0); -- 
    accessMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(16);
      gj_accessMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_update_start_
      -- CP-element group 15: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Update/$entry
      -- CP-element group 15: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_144_delayed_4_0_143_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(15), ack => W_read_write_bar_144_delayed_4_0_143_inst_req_1); -- 
    accessMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(17) & accessMem_CP_0_elements(20);
      gj_accessMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	2 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_sample_completed_
      -- CP-element group 16: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_144_delayed_4_0_143_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_144_delayed_4_0_143_inst_ack_0, ack => accessMem_CP_0_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_update_completed_
      -- CP-element group 17: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Update/$exit
      -- CP-element group 17: 	 assign_stmt_137_to_assign_stmt_151/assign_stmt_145_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_144_delayed_4_0_143_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_144_delayed_4_0_143_inst_ack_1, ack => accessMem_CP_0_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: 	9 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_sample_start_
      -- CP-element group 18: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_start/$entry
      -- CP-element group 18: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_start/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_150_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(18), ack => MUX_150_inst_req_0); -- 
    accessMem_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(17) & accessMem_CP_0_elements(9) & accessMem_CP_0_elements(20);
      gj_accessMem_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_update_start_
      -- CP-element group 19: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_complete/$entry
      -- CP-element group 19: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_complete/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_150_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(19), ack => MUX_150_inst_req_1); -- 
    accessMem_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(5) & accessMem_CP_0_elements(21);
      gj_accessMem_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	7 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_sample_completed_
      -- CP-element group 20: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_start/$exit
      -- CP-element group 20: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_start/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_150_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_150_inst_ack_0, ack => accessMem_CP_0_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_update_completed_
      -- CP-element group 21: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_complete/$exit
      -- CP-element group 21: 	 assign_stmt_137_to_assign_stmt_151/MUX_150_complete/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_150_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_150_inst_ack_1, ack => accessMem_CP_0_elements(21)); -- 
    -- CP-element group 22:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	10 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 assign_stmt_137_to_assign_stmt_151/array_obj_ref_136_array_obj_ref_140_delay
      -- 
    -- logger for CP element group accessMem_CP_0_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_CP_0_elements(22) is a control-delay.
    cp_element_22_delay: control_delay_element  generic map(name => " 22_delay", delay_value => 1)  port map(req => accessMem_CP_0_elements(8), ack => accessMem_CP_0_elements(22), clk => clk, reset =>reset);
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	12 
    -- CP-element group 23: 	13 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	28 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 assign_stmt_137_to_assign_stmt_151/$exit
      -- 
    -- logger for CP element group accessMem_CP_0_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(12) & accessMem_CP_0_elements(13) & accessMem_CP_0_elements(21);
      gj_accessMem_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  place  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 read_write_bar_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(24) <= accessMem_CP_0_elements(2);
    -- CP-element group 25:  place  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	3 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 addr_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(25) <= accessMem_CP_0_elements(3);
    -- CP-element group 26:  place  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	4 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 write_data_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(26) <= accessMem_CP_0_elements(4);
    -- CP-element group 27:  place  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	5 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 read_data_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 28:  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 $exit
      -- 
    -- logger for CP element group accessMem_CP_0_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(28) <= accessMem_CP_0_elements(23);
    --  hookup: inputs to control-path 
    accessMem_CP_0_elements(27) <= read_data_update_enable;
    -- hookup: output from control-path 
    read_write_bar_update_enable <= accessMem_CP_0_elements(24);
    addr_update_enable <= accessMem_CP_0_elements(25);
    write_data_update_enable <= accessMem_CP_0_elements(26);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_addr_135_resized : std_logic_vector(9 downto 0);
    signal R_addr_135_scaled : std_logic_vector(9 downto 0);
    signal R_addr_139_resized : std_logic_vector(9 downto 0);
    signal R_addr_139_scaled : std_logic_vector(9 downto 0);
    signal array_obj_ref_136_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_136_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_136_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_136_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_136_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_136_word_address_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_136_word_offset_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_140_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_140_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_140_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_140_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_140_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_140_word_address_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_140_word_offset_0 : std_logic_vector(9 downto 0);
    signal konst_149_wire_constant : std_logic_vector(31 downto 0);
    signal read_write_bar_144_delayed_4_0_145 : std_logic_vector(0 downto 0);
    signal t_read_data_137 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_136_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_136_resized_base_address <= "0000000000";
    array_obj_ref_136_word_offset_0 <= "0000000000";
    array_obj_ref_140_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_140_resized_base_address <= "0000000000";
    array_obj_ref_140_word_offset_0 <= "0000000000";
    konst_149_wire_constant <= "00000000000000000000000000000000";
    -- logger for split-operator MUX_150_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_150_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:MUX_150_inst:started:   inputs: " & " read_write_bar_144_delayed_4_0_145 = "& Convert_SLV_To_Hex_String(read_write_bar_144_delayed_4_0_145) & " t_read_data_137 = "& Convert_SLV_To_Hex_String(t_read_data_137) & " konst_149_wire_constant = "& Convert_SLV_To_Hex_String(konst_149_wire_constant));
          --
        end if; 
        if MUX_150_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:MUX_150_inst:finished:  outputs: " & " read_data_buffer= "  & Convert_SLV_To_Hex_String(read_data_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_150_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_150_inst_req_0;
      MUX_150_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_150_inst_req_1;
      MUX_150_inst_ack_1<= update_ack(0);
      MUX_150_inst: SelectSplitProtocol generic map(name => "MUX_150_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => t_read_data_137, y => konst_149_wire_constant, sel => read_write_bar_144_delayed_4_0_145, z => read_data_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator W_read_write_bar_144_delayed_4_0_143_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_144_delayed_4_0_143_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_144_delayed_4_0_143_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_144_delayed_4_0_143_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_144_delayed_4_0_143_inst:finished:  outputs: " & " read_write_bar_144_delayed_4_0_145= "  & Convert_SLV_To_Hex_String(read_write_bar_144_delayed_4_0_145));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_144_delayed_4_0_143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_144_delayed_4_0_143_inst_req_0;
      W_read_write_bar_144_delayed_4_0_143_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_144_delayed_4_0_143_inst_req_1;
      W_read_write_bar_144_delayed_4_0_143_inst_ack_1<= rack(0);
      W_read_write_bar_144_delayed_4_0_143_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_144_delayed_4_0_143_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_144_delayed_4_0_145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_136_addr_0 flow-through 
    process(array_obj_ref_136_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_addr_0:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_136_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_136_root_address) & "outputs: " & " array_obj_ref_136_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_136_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_136_addr_0
    process(array_obj_ref_136_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_136_root_address;
      ov(9 downto 0) := iv;
      array_obj_ref_136_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_136_gather_scatter flow-through 
    process(t_read_data_137) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_gather_scatter:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_136_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_136_data_0) & "outputs: " & " t_read_data_137= "  & Convert_SLV_To_Hex_String(t_read_data_137));
      --
    end process; 
    -- equivalence array_obj_ref_136_gather_scatter
    process(array_obj_ref_136_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_136_data_0;
      ov(31 downto 0) := iv;
      t_read_data_137 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_136_index_0_rename flow-through 
    process(R_addr_135_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_index_0_rename:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_135_resized = "& Convert_SLV_To_Hex_String(R_addr_135_resized) & "outputs: " & " R_addr_135_scaled= "  & Convert_SLV_To_Hex_String(R_addr_135_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_136_index_0_rename
    process(R_addr_135_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_135_resized;
      ov(9 downto 0) := iv;
      R_addr_135_scaled <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_136_index_0_resize flow-through 
    process(R_addr_135_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_index_0_resize:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_135_resized= "  & Convert_SLV_To_Hex_String(R_addr_135_resized));
      --
    end process; 
    -- equivalence array_obj_ref_136_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov(9 downto 0) := iv;
      R_addr_135_resized <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_136_index_offset flow-through 
    process(array_obj_ref_136_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_index_offset:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_135_scaled = "& Convert_SLV_To_Hex_String(R_addr_135_scaled) & "outputs: " & " array_obj_ref_136_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_136_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_136_index_offset
    process(R_addr_135_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_135_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_136_final_offset <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_136_root_address_inst flow-through 
    process(array_obj_ref_136_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_root_address_inst:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_136_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_136_final_offset) & "outputs: " & " array_obj_ref_136_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_136_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_136_root_address_inst
    process(array_obj_ref_136_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_136_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_136_root_address <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_140_addr_0 flow-through 
    process(array_obj_ref_140_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_addr_0:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_140_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_140_root_address) & "outputs: " & " array_obj_ref_140_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_140_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_140_addr_0
    process(array_obj_ref_140_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_140_root_address;
      ov(9 downto 0) := iv;
      array_obj_ref_140_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_140_gather_scatter flow-through 
    process(array_obj_ref_140_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_gather_scatter:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " write_data_buffer = "& Convert_SLV_To_Hex_String(write_data_buffer) & "outputs: " & " array_obj_ref_140_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_140_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_140_gather_scatter
    process(write_data_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := write_data_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_140_data_0 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_140_index_0_rename flow-through 
    process(R_addr_139_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_index_0_rename:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_139_resized = "& Convert_SLV_To_Hex_String(R_addr_139_resized) & "outputs: " & " R_addr_139_scaled= "  & Convert_SLV_To_Hex_String(R_addr_139_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_140_index_0_rename
    process(R_addr_139_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_139_resized;
      ov(9 downto 0) := iv;
      R_addr_139_scaled <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_140_index_0_resize flow-through 
    process(R_addr_139_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_index_0_resize:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_139_resized= "  & Convert_SLV_To_Hex_String(R_addr_139_resized));
      --
    end process; 
    -- equivalence array_obj_ref_140_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov(9 downto 0) := iv;
      R_addr_139_resized <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_140_index_offset flow-through 
    process(array_obj_ref_140_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_index_offset:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_139_scaled = "& Convert_SLV_To_Hex_String(R_addr_139_scaled) & "outputs: " & " array_obj_ref_140_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_140_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_140_index_offset
    process(R_addr_139_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_139_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_140_final_offset <= ov(9 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_140_root_address_inst flow-through 
    process(array_obj_ref_140_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_root_address_inst:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_140_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_140_final_offset) & "outputs: " & " array_obj_ref_140_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_140_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_140_root_address_inst
    process(array_obj_ref_140_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_140_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_140_root_address <= ov(9 downto 0);
      --
    end process;
    -- logger for split-operator array_obj_ref_136_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_136_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_load_0:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_136_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_136_word_address_0));
          --
        end if; 
        if array_obj_ref_136_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_136_load_0:finished:  outputs: " & " array_obj_ref_136_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_136_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_136_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_136_load_0_req_0,
        array_obj_ref_136_load_0_ack_0,
        array_obj_ref_136_load_0_req_1,
        array_obj_ref_136_load_0_ack_1,
        "array_obj_ref_136_load_0",
        "memory_space_0" ,
        array_obj_ref_136_data_0,
        array_obj_ref_136_word_address_0,
        "array_obj_ref_136_data_0",
        "array_obj_ref_136_word_address_0" -- 
      );
      reqL_unguarded(0) <= array_obj_ref_136_load_0_req_0;
      array_obj_ref_136_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_136_load_0_req_1;
      array_obj_ref_136_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_136_word_address_0;
      array_obj_ref_136_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 10,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(9 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator array_obj_ref_140_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_140_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_store_0:started:   inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_140_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_140_word_address_0) & " array_obj_ref_140_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_140_data_0));
          --
        end if; 
        if array_obj_ref_140_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_140_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_140_store_0_req_0,
      array_obj_ref_140_store_0_ack_0,
      array_obj_ref_140_store_0_req_1,
      array_obj_ref_140_store_0_ack_1,
      "array_obj_ref_140_store_0",
      "memory_space_0" ,
      array_obj_ref_140_data_0,
      array_obj_ref_140_word_address_0,
      "array_obj_ref_140_data_0",
      "array_obj_ref_140_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_140_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_140_store_0_req_0;
      array_obj_ref_140_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_140_store_0_req_1;
      array_obj_ref_140_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_140_word_address_0;
      data_in <= array_obj_ref_140_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(9 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessReg is -- 
  generic (tag_length : integer); 
  port ( -- 
    valid_1 : in  std_logic_vector(0 downto 0);
    addr_1 : in  std_logic_vector(7 downto 0);
    valid_2 : in  std_logic_vector(0 downto 0);
    addr_2 : in  std_logic_vector(7 downto 0);
    valid_w : in  std_logic_vector(0 downto 0);
    addr_w : in  std_logic_vector(7 downto 0);
    data_to_be_written : in  std_logic_vector(31 downto 0);
    read_data_1 : out  std_logic_vector(31 downto 0);
    read_data_2 : out  std_logic_vector(31 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessReg;
architecture accessReg_arch of accessReg is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 59)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal valid_1_buffer :  std_logic_vector(0 downto 0);
  signal valid_1_update_enable: Boolean;
  signal addr_1_buffer :  std_logic_vector(7 downto 0);
  signal addr_1_update_enable: Boolean;
  signal valid_2_buffer :  std_logic_vector(0 downto 0);
  signal valid_2_update_enable: Boolean;
  signal addr_2_buffer :  std_logic_vector(7 downto 0);
  signal addr_2_update_enable: Boolean;
  signal valid_w_buffer :  std_logic_vector(0 downto 0);
  signal valid_w_update_enable: Boolean;
  signal addr_w_buffer :  std_logic_vector(7 downto 0);
  signal addr_w_update_enable: Boolean;
  signal data_to_be_written_buffer :  std_logic_vector(31 downto 0);
  signal data_to_be_written_update_enable: Boolean;
  -- output port buffer signals
  signal read_data_1_buffer :  std_logic_vector(31 downto 0);
  signal read_data_1_update_enable: Boolean;
  signal read_data_2_buffer :  std_logic_vector(31 downto 0);
  signal read_data_2_update_enable: Boolean;
  signal accessReg_CP_173_start: Boolean;
  signal accessReg_CP_173_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_166_load_0_req_0 : boolean;
  signal array_obj_ref_166_load_0_ack_0 : boolean;
  signal array_obj_ref_166_load_0_req_1 : boolean;
  signal array_obj_ref_166_load_0_ack_1 : boolean;
  signal array_obj_ref_171_load_0_req_0 : boolean;
  signal array_obj_ref_171_load_0_ack_0 : boolean;
  signal array_obj_ref_171_load_0_req_1 : boolean;
  signal array_obj_ref_171_load_0_ack_1 : boolean;
  signal W_valid_1_171_delayed_4_0_173_inst_req_0 : boolean;
  signal W_valid_1_171_delayed_4_0_173_inst_ack_0 : boolean;
  signal W_valid_1_171_delayed_4_0_173_inst_req_1 : boolean;
  signal W_valid_1_171_delayed_4_0_173_inst_ack_1 : boolean;
  signal MUX_180_inst_req_0 : boolean;
  signal MUX_180_inst_ack_0 : boolean;
  signal MUX_180_inst_req_1 : boolean;
  signal MUX_180_inst_ack_1 : boolean;
  signal W_valid_2_177_delayed_4_0_182_inst_req_0 : boolean;
  signal W_valid_2_177_delayed_4_0_182_inst_ack_0 : boolean;
  signal W_valid_2_177_delayed_4_0_182_inst_req_1 : boolean;
  signal W_valid_2_177_delayed_4_0_182_inst_ack_1 : boolean;
  signal MUX_189_inst_req_0 : boolean;
  signal MUX_189_inst_ack_0 : boolean;
  signal MUX_189_inst_req_1 : boolean;
  signal MUX_189_inst_ack_1 : boolean;
  signal array_obj_ref_193_store_0_req_0 : boolean;
  signal array_obj_ref_193_store_0_ack_0 : boolean;
  signal array_obj_ref_193_store_0_req_1 : boolean;
  signal array_obj_ref_193_store_0_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessReg_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 59) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= valid_1;
  valid_1_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(8 downto 1) <= addr_1;
  addr_1_buffer <= in_buffer_data_out(8 downto 1);
  in_buffer_data_in(9 downto 9) <= valid_2;
  valid_2_buffer <= in_buffer_data_out(9 downto 9);
  in_buffer_data_in(17 downto 10) <= addr_2;
  addr_2_buffer <= in_buffer_data_out(17 downto 10);
  in_buffer_data_in(18 downto 18) <= valid_w;
  valid_w_buffer <= in_buffer_data_out(18 downto 18);
  in_buffer_data_in(26 downto 19) <= addr_w;
  addr_w_buffer <= in_buffer_data_out(26 downto 19);
  in_buffer_data_in(58 downto 27) <= data_to_be_written;
  data_to_be_written_buffer <= in_buffer_data_out(58 downto 27);
  in_buffer_data_in(tag_length + 58 downto 59) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 58 downto 59);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 8) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1,8 => 7);
    constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1,8 => 7);
    constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 9); -- 
  begin -- 
    preds <= valid_1_update_enable & addr_1_update_enable & valid_2_update_enable & addr_2_update_enable & valid_w_update_enable & addr_w_update_enable & data_to_be_written_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessReg_CP_173_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessReg_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= read_data_1_buffer;
  read_data_1 <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= read_data_2_buffer;
  read_data_2 <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessReg_CP_173_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  read_data_1_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "read_data_1_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_data_1_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_data_1_update_enable, clk => clk, reset => reset); --
  end block;
  read_data_2_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "read_data_2_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_data_2_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_data_2_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessReg_CP_173_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessReg_CP_173_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accessReg_CP_173_start,"accessReg cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accessReg_CP_173_symbol, "accessReg cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessReg_CP_173: Block -- control-path 
    signal accessReg_CP_173_elements: BooleanArray(51 downto 0);
    -- 
  begin -- 
    accessReg_CP_173_elements(0) <= accessReg_CP_173_start;
    accessReg_CP_173_symbol <= accessReg_CP_173_elements(51);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group accessReg_CP_173_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	15 
    -- CP-element group 1: 	19 
    -- CP-element group 1: 	27 
    -- CP-element group 1: 	35 
    -- CP-element group 1: 	11 
    -- CP-element group 1:  members (79) 
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_offset_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_resized_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_computed_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_word_addrgen/root_register_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_offset_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_resized_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_computed_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_word_addrgen/root_register_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_offset_calculated
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_resized_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_computed_0
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(1) <= accessReg_CP_173_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	13 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	42 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_195/valid_1_update_enable
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_195/valid_1_update_enable_out
      -- 
    -- logger for CP element group accessReg_CP_173_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessReg_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(21) & accessReg_CP_173_elements(13);
      gj_accessReg_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	13 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	43 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_195/addr_1_update_enable
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_195/addr_1_update_enable_out
      -- 
    -- logger for CP element group accessReg_CP_173_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessReg_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessReg_CP_173_elements(13);
      gj_accessReg_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	17 
    -- CP-element group 4: 	29 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	44 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_167_to_assign_stmt_195/valid_2_update_enable
      -- CP-element group 4: 	 assign_stmt_167_to_assign_stmt_195/valid_2_update_enable_out
      -- 
    -- logger for CP element group accessReg_CP_173_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessReg_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(17) & accessReg_CP_173_elements(29);
      gj_accessReg_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	17 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	45 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_195/addr_2_update_enable
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_195/addr_2_update_enable_out
      -- 
    -- logger for CP element group accessReg_CP_173_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessReg_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessReg_CP_173_elements(17);
      gj_accessReg_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	37 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	46 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_167_to_assign_stmt_195/valid_w_update_enable
      -- CP-element group 6: 	 assign_stmt_167_to_assign_stmt_195/valid_w_update_enable_out
      -- 
    -- logger for CP element group accessReg_CP_173_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessReg_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessReg_CP_173_elements(37);
      gj_accessReg_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	37 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	47 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_167_to_assign_stmt_195/addr_w_update_enable
      -- CP-element group 7: 	 assign_stmt_167_to_assign_stmt_195/addr_w_update_enable_out
      -- 
    -- logger for CP element group accessReg_CP_173_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessReg_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessReg_CP_173_elements(37);
      gj_accessReg_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	37 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	48 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 assign_stmt_167_to_assign_stmt_195/data_to_be_written_update_enable
      -- CP-element group 8: 	 assign_stmt_167_to_assign_stmt_195/data_to_be_written_update_enable_out
      -- 
    -- logger for CP element group accessReg_CP_173_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessReg_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessReg_CP_173_elements(37);
      gj_accessReg_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	49 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	24 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 assign_stmt_167_to_assign_stmt_195/read_data_1_update_enable
      -- CP-element group 9: 	 assign_stmt_167_to_assign_stmt_195/read_data_1_update_enable_in
      -- 
    -- logger for CP element group accessReg_CP_173_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(9) <= accessReg_CP_173_elements(49);
    -- CP-element group 10:  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	50 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	32 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 assign_stmt_167_to_assign_stmt_195/read_data_2_update_enable
      -- CP-element group 10: 	 assign_stmt_167_to_assign_stmt_195/read_data_2_update_enable_in
      -- 
    -- logger for CP element group accessReg_CP_173_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(10) <= accessReg_CP_173_elements(50);
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_sample_start_
      -- CP-element group 11: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/word_access_start/$entry
      -- CP-element group 11: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/word_access_start/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessReg_CP_173_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_166_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(11), ack => array_obj_ref_166_load_0_req_0); -- 
    accessReg_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(1) & accessReg_CP_173_elements(37) & accessReg_CP_173_elements(13);
      gj_accessReg_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	25 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_update_start_
      -- CP-element group 12: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/$entry
      -- CP-element group 12: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/word_access_complete/$entry
      -- CP-element group 12: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/word_access_complete/word_0/$entry
      -- CP-element group 12: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessReg_CP_173_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_166_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(12), ack => array_obj_ref_166_load_0_req_1); -- 
    accessReg_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(14) & accessReg_CP_173_elements(25);
      gj_accessReg_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	39 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: 	11 
    -- CP-element group 13: 	3 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_sample_completed_
      -- CP-element group 13: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/word_access_start/$exit
      -- CP-element group 13: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessReg_CP_173_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_166_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_166_load_0_ack_0, ack => accessReg_CP_173_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	23 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_update_completed_
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/$exit
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/word_access_complete/$exit
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/array_obj_ref_166_Merge/$entry
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/array_obj_ref_166_Merge/$exit
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/array_obj_ref_166_Merge/merge_req
      -- CP-element group 14: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_Update/array_obj_ref_166_Merge/merge_ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_166_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_166_load_0_ack_1, ack => accessReg_CP_173_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	1 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	37 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_sample_start_
      -- CP-element group 15: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/$entry
      -- CP-element group 15: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/word_access_start/$entry
      -- CP-element group 15: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessReg_CP_173_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_171_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(15), ack => array_obj_ref_171_load_0_req_0); -- 
    accessReg_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(1) & accessReg_CP_173_elements(17) & accessReg_CP_173_elements(37);
      gj_accessReg_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	33 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_update_start_
      -- CP-element group 16: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/$entry
      -- CP-element group 16: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/word_access_complete/$entry
      -- CP-element group 16: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/word_access_complete/word_0/$entry
      -- CP-element group 16: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessReg_CP_173_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_171_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(16), ack => array_obj_ref_171_load_0_req_1); -- 
    accessReg_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(18) & accessReg_CP_173_elements(33);
      gj_accessReg_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	40 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: 	5 
    -- CP-element group 17: 	4 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_sample_completed_
      -- CP-element group 17: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/$exit
      -- CP-element group 17: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/word_access_start/$exit
      -- CP-element group 17: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessReg_CP_173_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_171_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_171_load_0_ack_0, ack => accessReg_CP_173_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	31 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_update_completed_
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/$exit
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/word_access_complete/$exit
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/array_obj_ref_171_Merge/$entry
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/array_obj_ref_171_Merge/$exit
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/array_obj_ref_171_Merge/merge_req
      -- CP-element group 18: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_Update/array_obj_ref_171_Merge/merge_ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_171_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_171_load_0_ack_1, ack => accessReg_CP_173_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	1 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_sample_start_
      -- CP-element group 19: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Sample/$entry
      -- CP-element group 19: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Sample/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_1_171_delayed_4_0_173_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(19), ack => W_valid_1_171_delayed_4_0_173_inst_req_0); -- 
    accessReg_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(1) & accessReg_CP_173_elements(21);
      gj_accessReg_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: 	25 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_update_start_
      -- CP-element group 20: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Update/$entry
      -- CP-element group 20: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Update/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_1_171_delayed_4_0_173_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(20), ack => W_valid_1_171_delayed_4_0_173_inst_req_1); -- 
    accessReg_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(22) & accessReg_CP_173_elements(25);
      gj_accessReg_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: 	2 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_sample_completed_
      -- CP-element group 21: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Sample/$exit
      -- CP-element group 21: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Sample/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_1_171_delayed_4_0_173_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_valid_1_171_delayed_4_0_173_inst_ack_0, ack => accessReg_CP_173_elements(21)); -- 
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	20 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_update_completed_
      -- CP-element group 22: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Update/$exit
      -- CP-element group 22: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_175_Update/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_1_171_delayed_4_0_173_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_valid_1_171_delayed_4_0_173_inst_ack_1, ack => accessReg_CP_173_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	14 
    -- CP-element group 23: 	22 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_sample_start_
      -- CP-element group 23: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_start/$entry
      -- CP-element group 23: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_start/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_180_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(23), ack => MUX_180_inst_req_0); -- 
    accessReg_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(14) & accessReg_CP_173_elements(22) & accessReg_CP_173_elements(25);
      gj_accessReg_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	9 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_update_start_
      -- CP-element group 24: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_complete/$entry
      -- CP-element group 24: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_complete/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_180_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(24), ack => MUX_180_inst_req_1); -- 
    accessReg_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(9) & accessReg_CP_173_elements(26);
      gj_accessReg_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	23 
    -- CP-element group 25: 	12 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_sample_completed_
      -- CP-element group 25: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_start/$exit
      -- CP-element group 25: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_start/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_180_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_180_inst_ack_0, ack => accessReg_CP_173_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	41 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_update_completed_
      -- CP-element group 26: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_complete/$exit
      -- CP-element group 26: 	 assign_stmt_167_to_assign_stmt_195/MUX_180_complete/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_180_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_180_inst_ack_1, ack => accessReg_CP_173_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	1 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_sample_start_
      -- CP-element group 27: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Sample/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_2_177_delayed_4_0_182_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(27), ack => W_valid_2_177_delayed_4_0_182_inst_req_0); -- 
    accessReg_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(1) & accessReg_CP_173_elements(29);
      gj_accessReg_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: 	33 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_update_start_
      -- CP-element group 28: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Update/$entry
      -- CP-element group 28: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Update/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_2_177_delayed_4_0_182_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(28), ack => W_valid_2_177_delayed_4_0_182_inst_req_1); -- 
    accessReg_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(30) & accessReg_CP_173_elements(33);
      gj_accessReg_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: 	4 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_sample_completed_
      -- CP-element group 29: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Sample/$exit
      -- CP-element group 29: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Sample/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_2_177_delayed_4_0_182_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_valid_2_177_delayed_4_0_182_inst_ack_0, ack => accessReg_CP_173_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_update_completed_
      -- CP-element group 30: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Update/$exit
      -- CP-element group 30: 	 assign_stmt_167_to_assign_stmt_195/assign_stmt_184_Update/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:W_valid_2_177_delayed_4_0_182_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_valid_2_177_delayed_4_0_182_inst_ack_1, ack => accessReg_CP_173_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	30 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_sample_start_
      -- CP-element group 31: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_start/$entry
      -- CP-element group 31: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_start/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_189_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(31), ack => MUX_189_inst_req_0); -- 
    accessReg_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(18) & accessReg_CP_173_elements(30) & accessReg_CP_173_elements(33);
      gj_accessReg_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	10 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_update_start_
      -- CP-element group 32: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_complete/$entry
      -- CP-element group 32: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_complete/req
      -- 
    -- logger for CP element group accessReg_CP_173_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_189_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(32), ack => MUX_189_inst_req_1); -- 
    accessReg_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(10) & accessReg_CP_173_elements(34);
      gj_accessReg_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_sample_completed_
      -- CP-element group 33: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_start/$exit
      -- CP-element group 33: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_start/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_189_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_189_inst_ack_0, ack => accessReg_CP_173_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	41 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_update_completed_
      -- CP-element group 34: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_complete/$exit
      -- CP-element group 34: 	 assign_stmt_167_to_assign_stmt_195/MUX_189_complete/ack
      -- 
    -- logger for CP element group accessReg_CP_173_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:MUX_189_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_189_inst_ack_1, ack => accessReg_CP_173_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	1 
    -- CP-element group 35: 	39 
    -- CP-element group 35: 	40 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_sample_start_
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/$entry
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/array_obj_ref_193_Split/$entry
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/array_obj_ref_193_Split/$exit
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/array_obj_ref_193_Split/split_req
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/array_obj_ref_193_Split/split_ack
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/word_access_start/$entry
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/word_access_start/word_0/$entry
      -- CP-element group 35: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessReg_CP_173_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_193_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(35), ack => array_obj_ref_193_store_0_req_0); -- 
    accessReg_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(1) & accessReg_CP_173_elements(39) & accessReg_CP_173_elements(40) & accessReg_CP_173_elements(37);
      gj_accessReg_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_update_start_
      -- CP-element group 36: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/$entry
      -- CP-element group 36: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/word_access_complete/$entry
      -- CP-element group 36: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/word_access_complete/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessReg_CP_173_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_193_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessReg_CP_173_elements(36), ack => array_obj_ref_193_store_0_req_1); -- 
    accessReg_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessReg_CP_173_elements(38);
      gj_accessReg_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	41 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	15 
    -- CP-element group 37: 	35 
    -- CP-element group 37: 	11 
    -- CP-element group 37: 	8 
    -- CP-element group 37: 	7 
    -- CP-element group 37: 	6 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_sample_completed_
      -- CP-element group 37: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/$exit
      -- CP-element group 37: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/word_access_start/$exit
      -- CP-element group 37: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Sample/word_access_start/word_0/ra
      -- CP-element group 37: 	 assign_stmt_167_to_assign_stmt_195/ring_reenable_memory_space_1
      -- 
    -- logger for CP element group accessReg_CP_173_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_193_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_193_store_0_ack_0, ack => accessReg_CP_173_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_update_completed_
      -- CP-element group 38: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/$exit
      -- CP-element group 38: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/word_access_complete/$exit
      -- CP-element group 38: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/word_access_complete/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_193_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group accessReg_CP_173_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:array_obj_ref_193_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_193_store_0_ack_1, ack => accessReg_CP_173_elements(38)); -- 
    -- CP-element group 39:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	13 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	35 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_166_array_obj_ref_193_delay
      -- 
    -- logger for CP element group accessReg_CP_173_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessReg_CP_173_elements(39) is a control-delay.
    cp_element_39_delay: control_delay_element  generic map(name => " 39_delay", delay_value => 1)  port map(req => accessReg_CP_173_elements(13), ack => accessReg_CP_173_elements(39), clk => clk, reset =>reset);
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	35 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 assign_stmt_167_to_assign_stmt_195/array_obj_ref_171_array_obj_ref_193_delay
      -- 
    -- logger for CP element group accessReg_CP_173_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessReg_CP_173_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => accessReg_CP_173_elements(17), ack => accessReg_CP_173_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	26 
    -- CP-element group 41: 	34 
    -- CP-element group 41: 	37 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	51 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 assign_stmt_167_to_assign_stmt_195/$exit
      -- 
    -- logger for CP element group accessReg_CP_173_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "accessReg_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessReg_CP_173_elements(26) & accessReg_CP_173_elements(34) & accessReg_CP_173_elements(37) & accessReg_CP_173_elements(38);
      gj_accessReg_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessReg_CP_173_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  place  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	2 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 valid_1_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(42) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(42) <= accessReg_CP_173_elements(2);
    -- CP-element group 43:  place  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	3 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 addr_1_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(43) <= accessReg_CP_173_elements(3);
    -- CP-element group 44:  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	4 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 valid_2_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(44) <= accessReg_CP_173_elements(4);
    -- CP-element group 45:  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	5 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 addr_2_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(45) <= accessReg_CP_173_elements(5);
    -- CP-element group 46:  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	6 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 valid_w_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(46) <= accessReg_CP_173_elements(6);
    -- CP-element group 47:  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	7 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 addr_w_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(47) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(47) <= accessReg_CP_173_elements(7);
    -- CP-element group 48:  place  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	8 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 data_to_be_written_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(48) <= accessReg_CP_173_elements(8);
    -- CP-element group 49:  place  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	9 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 read_data_1_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 50:  place  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	10 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 read_data_2_update_enable
      -- 
    -- logger for CP element group accessReg_CP_173_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(50) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 51:  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	41 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 $exit
      -- 
    -- logger for CP element group accessReg_CP_173_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessReg_CP_173_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessReg:CP:accessReg_CP_173_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    accessReg_CP_173_elements(51) <= accessReg_CP_173_elements(41);
    --  hookup: inputs to control-path 
    accessReg_CP_173_elements(49) <= read_data_1_update_enable;
    accessReg_CP_173_elements(50) <= read_data_2_update_enable;
    -- hookup: output from control-path 
    valid_1_update_enable <= accessReg_CP_173_elements(42);
    addr_1_update_enable <= accessReg_CP_173_elements(43);
    valid_2_update_enable <= accessReg_CP_173_elements(44);
    addr_2_update_enable <= accessReg_CP_173_elements(45);
    valid_w_update_enable <= accessReg_CP_173_elements(46);
    addr_w_update_enable <= accessReg_CP_173_elements(47);
    data_to_be_written_update_enable <= accessReg_CP_173_elements(48);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_addr_1_165_resized : std_logic_vector(5 downto 0);
    signal R_addr_1_165_scaled : std_logic_vector(5 downto 0);
    signal R_addr_2_170_resized : std_logic_vector(5 downto 0);
    signal R_addr_2_170_scaled : std_logic_vector(5 downto 0);
    signal R_addr_w_192_resized : std_logic_vector(5 downto 0);
    signal R_addr_w_192_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_166_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_166_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_166_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_166_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_166_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_166_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_166_word_offset_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_171_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_171_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_171_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_171_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_171_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_171_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_171_word_offset_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_193_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_word_offset_0 : std_logic_vector(5 downto 0);
    signal konst_179_wire_constant : std_logic_vector(31 downto 0);
    signal konst_188_wire_constant : std_logic_vector(31 downto 0);
    signal t_read_data_1_167 : std_logic_vector(31 downto 0);
    signal t_read_data_2_172 : std_logic_vector(31 downto 0);
    signal valid_1_171_delayed_4_0_175 : std_logic_vector(0 downto 0);
    signal valid_2_177_delayed_4_0_184 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_166_offset_scale_factor_0 <= "000001";
    array_obj_ref_166_resized_base_address <= "000000";
    array_obj_ref_166_word_offset_0 <= "000000";
    array_obj_ref_171_offset_scale_factor_0 <= "000001";
    array_obj_ref_171_resized_base_address <= "000000";
    array_obj_ref_171_word_offset_0 <= "000000";
    array_obj_ref_193_offset_scale_factor_0 <= "000001";
    array_obj_ref_193_resized_base_address <= "000000";
    array_obj_ref_193_word_offset_0 <= "000000";
    konst_179_wire_constant <= "00000000000000000000000000000000";
    konst_188_wire_constant <= "00000000000000000000000000000000";
    -- logger for split-operator MUX_180_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_180_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:MUX_180_inst:started:   inputs: " & " valid_1_171_delayed_4_0_175 = "& Convert_SLV_To_Hex_String(valid_1_171_delayed_4_0_175) & " t_read_data_1_167 = "& Convert_SLV_To_Hex_String(t_read_data_1_167) & " konst_179_wire_constant = "& Convert_SLV_To_Hex_String(konst_179_wire_constant));
          --
        end if; 
        if MUX_180_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:MUX_180_inst:finished:  outputs: " & " read_data_1_buffer= "  & Convert_SLV_To_Hex_String(read_data_1_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_180_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_180_inst_req_0;
      MUX_180_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_180_inst_req_1;
      MUX_180_inst_ack_1<= update_ack(0);
      MUX_180_inst: SelectSplitProtocol generic map(name => "MUX_180_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => t_read_data_1_167, y => konst_179_wire_constant, sel => valid_1_171_delayed_4_0_175, z => read_data_1_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator MUX_189_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_189_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:MUX_189_inst:started:   inputs: " & " valid_2_177_delayed_4_0_184 = "& Convert_SLV_To_Hex_String(valid_2_177_delayed_4_0_184) & " t_read_data_2_172 = "& Convert_SLV_To_Hex_String(t_read_data_2_172) & " konst_188_wire_constant = "& Convert_SLV_To_Hex_String(konst_188_wire_constant));
          --
        end if; 
        if MUX_189_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:MUX_189_inst:finished:  outputs: " & " read_data_2_buffer= "  & Convert_SLV_To_Hex_String(read_data_2_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_189_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_189_inst_req_0;
      MUX_189_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_189_inst_req_1;
      MUX_189_inst_ack_1<= update_ack(0);
      MUX_189_inst: SelectSplitProtocol generic map(name => "MUX_189_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => t_read_data_2_172, y => konst_188_wire_constant, sel => valid_2_177_delayed_4_0_184, z => read_data_2_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator W_valid_1_171_delayed_4_0_173_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_valid_1_171_delayed_4_0_173_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:W_valid_1_171_delayed_4_0_173_inst:started:   inputs: " & " valid_1_buffer = "& Convert_SLV_To_Hex_String(valid_1_buffer));
          --
        end if; 
        if W_valid_1_171_delayed_4_0_173_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:W_valid_1_171_delayed_4_0_173_inst:finished:  outputs: " & " valid_1_171_delayed_4_0_175= "  & Convert_SLV_To_Hex_String(valid_1_171_delayed_4_0_175));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_valid_1_171_delayed_4_0_173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_valid_1_171_delayed_4_0_173_inst_req_0;
      W_valid_1_171_delayed_4_0_173_inst_ack_0<= wack(0);
      rreq(0) <= W_valid_1_171_delayed_4_0_173_inst_req_1;
      W_valid_1_171_delayed_4_0_173_inst_ack_1<= rack(0);
      W_valid_1_171_delayed_4_0_173_inst : InterlockBuffer generic map ( -- 
        name => "W_valid_1_171_delayed_4_0_173_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valid_1_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => valid_1_171_delayed_4_0_175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_valid_2_177_delayed_4_0_182_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_valid_2_177_delayed_4_0_182_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:W_valid_2_177_delayed_4_0_182_inst:started:   inputs: " & " valid_2_buffer = "& Convert_SLV_To_Hex_String(valid_2_buffer));
          --
        end if; 
        if W_valid_2_177_delayed_4_0_182_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:W_valid_2_177_delayed_4_0_182_inst:finished:  outputs: " & " valid_2_177_delayed_4_0_184= "  & Convert_SLV_To_Hex_String(valid_2_177_delayed_4_0_184));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_valid_2_177_delayed_4_0_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_valid_2_177_delayed_4_0_182_inst_req_0;
      W_valid_2_177_delayed_4_0_182_inst_ack_0<= wack(0);
      rreq(0) <= W_valid_2_177_delayed_4_0_182_inst_req_1;
      W_valid_2_177_delayed_4_0_182_inst_ack_1<= rack(0);
      W_valid_2_177_delayed_4_0_182_inst : InterlockBuffer generic map ( -- 
        name => "W_valid_2_177_delayed_4_0_182_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valid_2_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => valid_2_177_delayed_4_0_184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_166_addr_0 flow-through 
    process(array_obj_ref_166_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_addr_0:flowthrough  inputs: " & " valid_1_buffer (guard)= " & Convert_SLV_To_String(valid_1_buffer) & " array_obj_ref_166_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_166_root_address) & "outputs: " & " array_obj_ref_166_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_166_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_166_addr_0
    process(array_obj_ref_166_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_166_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_166_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_166_gather_scatter flow-through 
    process(t_read_data_1_167) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_gather_scatter:flowthrough  inputs: " & " valid_1_buffer (guard)= " & Convert_SLV_To_String(valid_1_buffer) & " array_obj_ref_166_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_166_data_0) & "outputs: " & " t_read_data_1_167= "  & Convert_SLV_To_Hex_String(t_read_data_1_167));
      --
    end process; 
    -- equivalence array_obj_ref_166_gather_scatter
    process(array_obj_ref_166_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_166_data_0;
      ov(31 downto 0) := iv;
      t_read_data_1_167 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_166_index_0_rename flow-through 
    process(R_addr_1_165_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_index_0_rename:flowthrough  inputs: " & " valid_1_buffer (guard)= " & Convert_SLV_To_String(valid_1_buffer) & " R_addr_1_165_resized = "& Convert_SLV_To_Hex_String(R_addr_1_165_resized) & "outputs: " & " R_addr_1_165_scaled= "  & Convert_SLV_To_Hex_String(R_addr_1_165_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_166_index_0_rename
    process(R_addr_1_165_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_1_165_resized;
      ov(5 downto 0) := iv;
      R_addr_1_165_scaled <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_166_index_0_resize flow-through 
    process(R_addr_1_165_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_index_0_resize:flowthrough  inputs: " & " valid_1_buffer (guard)= " & Convert_SLV_To_String(valid_1_buffer) & " addr_1_buffer = "& Convert_SLV_To_Hex_String(addr_1_buffer) & "outputs: " & " R_addr_1_165_resized= "  & Convert_SLV_To_Hex_String(R_addr_1_165_resized));
      --
    end process; 
    -- equivalence array_obj_ref_166_index_0_resize
    process(addr_1_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_1_buffer;
      ov := iv(5 downto 0);
      R_addr_1_165_resized <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_166_index_offset flow-through 
    process(array_obj_ref_166_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_index_offset:flowthrough  inputs: " & " valid_1_buffer (guard)= " & Convert_SLV_To_String(valid_1_buffer) & " R_addr_1_165_scaled = "& Convert_SLV_To_Hex_String(R_addr_1_165_scaled) & "outputs: " & " array_obj_ref_166_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_166_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_166_index_offset
    process(R_addr_1_165_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_1_165_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_166_final_offset <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_166_root_address_inst flow-through 
    process(array_obj_ref_166_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_root_address_inst:flowthrough  inputs: " & " valid_1_buffer (guard)= " & Convert_SLV_To_String(valid_1_buffer) & " array_obj_ref_166_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_166_final_offset) & "outputs: " & " array_obj_ref_166_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_166_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_166_root_address_inst
    process(array_obj_ref_166_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_166_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_166_root_address <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_171_addr_0 flow-through 
    process(array_obj_ref_171_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_addr_0:flowthrough  inputs: " & " valid_2_buffer (guard)= " & Convert_SLV_To_String(valid_2_buffer) & " array_obj_ref_171_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_171_root_address) & "outputs: " & " array_obj_ref_171_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_171_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_171_addr_0
    process(array_obj_ref_171_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_171_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_171_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_171_gather_scatter flow-through 
    process(t_read_data_2_172) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_gather_scatter:flowthrough  inputs: " & " valid_2_buffer (guard)= " & Convert_SLV_To_String(valid_2_buffer) & " array_obj_ref_171_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_171_data_0) & "outputs: " & " t_read_data_2_172= "  & Convert_SLV_To_Hex_String(t_read_data_2_172));
      --
    end process; 
    -- equivalence array_obj_ref_171_gather_scatter
    process(array_obj_ref_171_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_171_data_0;
      ov(31 downto 0) := iv;
      t_read_data_2_172 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_171_index_0_rename flow-through 
    process(R_addr_2_170_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_index_0_rename:flowthrough  inputs: " & " valid_2_buffer (guard)= " & Convert_SLV_To_String(valid_2_buffer) & " R_addr_2_170_resized = "& Convert_SLV_To_Hex_String(R_addr_2_170_resized) & "outputs: " & " R_addr_2_170_scaled= "  & Convert_SLV_To_Hex_String(R_addr_2_170_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_171_index_0_rename
    process(R_addr_2_170_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_2_170_resized;
      ov(5 downto 0) := iv;
      R_addr_2_170_scaled <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_171_index_0_resize flow-through 
    process(R_addr_2_170_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_index_0_resize:flowthrough  inputs: " & " valid_2_buffer (guard)= " & Convert_SLV_To_String(valid_2_buffer) & " addr_2_buffer = "& Convert_SLV_To_Hex_String(addr_2_buffer) & "outputs: " & " R_addr_2_170_resized= "  & Convert_SLV_To_Hex_String(R_addr_2_170_resized));
      --
    end process; 
    -- equivalence array_obj_ref_171_index_0_resize
    process(addr_2_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_2_buffer;
      ov := iv(5 downto 0);
      R_addr_2_170_resized <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_171_index_offset flow-through 
    process(array_obj_ref_171_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_index_offset:flowthrough  inputs: " & " valid_2_buffer (guard)= " & Convert_SLV_To_String(valid_2_buffer) & " R_addr_2_170_scaled = "& Convert_SLV_To_Hex_String(R_addr_2_170_scaled) & "outputs: " & " array_obj_ref_171_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_171_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_171_index_offset
    process(R_addr_2_170_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_2_170_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_171_final_offset <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_171_root_address_inst flow-through 
    process(array_obj_ref_171_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_root_address_inst:flowthrough  inputs: " & " valid_2_buffer (guard)= " & Convert_SLV_To_String(valid_2_buffer) & " array_obj_ref_171_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_171_final_offset) & "outputs: " & " array_obj_ref_171_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_171_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_171_root_address_inst
    process(array_obj_ref_171_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_171_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_171_root_address <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_addr_0 flow-through 
    process(array_obj_ref_193_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_addr_0:flowthrough  inputs: " & " valid_w_buffer (guard)= " & Convert_SLV_To_String(valid_w_buffer) & " array_obj_ref_193_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_193_root_address) & "outputs: " & " array_obj_ref_193_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_193_addr_0
    process(array_obj_ref_193_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_193_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_193_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_gather_scatter flow-through 
    process(array_obj_ref_193_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_gather_scatter:flowthrough  inputs: " & " valid_w_buffer (guard)= " & Convert_SLV_To_String(valid_w_buffer) & " data_to_be_written_buffer = "& Convert_SLV_To_Hex_String(data_to_be_written_buffer) & "outputs: " & " array_obj_ref_193_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_193_gather_scatter
    process(data_to_be_written_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := data_to_be_written_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_193_data_0 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_index_0_rename flow-through 
    process(R_addr_w_192_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_index_0_rename:flowthrough  inputs: " & " valid_w_buffer (guard)= " & Convert_SLV_To_String(valid_w_buffer) & " R_addr_w_192_resized = "& Convert_SLV_To_Hex_String(R_addr_w_192_resized) & "outputs: " & " R_addr_w_192_scaled= "  & Convert_SLV_To_Hex_String(R_addr_w_192_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_193_index_0_rename
    process(R_addr_w_192_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_w_192_resized;
      ov(5 downto 0) := iv;
      R_addr_w_192_scaled <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_index_0_resize flow-through 
    process(R_addr_w_192_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_index_0_resize:flowthrough  inputs: " & " valid_w_buffer (guard)= " & Convert_SLV_To_String(valid_w_buffer) & " addr_w_buffer = "& Convert_SLV_To_Hex_String(addr_w_buffer) & "outputs: " & " R_addr_w_192_resized= "  & Convert_SLV_To_Hex_String(R_addr_w_192_resized));
      --
    end process; 
    -- equivalence array_obj_ref_193_index_0_resize
    process(addr_w_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_w_buffer;
      ov := iv(5 downto 0);
      R_addr_w_192_resized <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_index_offset flow-through 
    process(array_obj_ref_193_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_index_offset:flowthrough  inputs: " & " valid_w_buffer (guard)= " & Convert_SLV_To_String(valid_w_buffer) & " R_addr_w_192_scaled = "& Convert_SLV_To_Hex_String(R_addr_w_192_scaled) & "outputs: " & " array_obj_ref_193_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_193_index_offset
    process(R_addr_w_192_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_w_192_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_193_final_offset <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_root_address_inst flow-through 
    process(array_obj_ref_193_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_root_address_inst:flowthrough  inputs: " & " valid_w_buffer (guard)= " & Convert_SLV_To_String(valid_w_buffer) & " array_obj_ref_193_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_193_final_offset) & "outputs: " & " array_obj_ref_193_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_193_root_address_inst
    process(array_obj_ref_193_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_193_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_193_root_address <= ov(5 downto 0);
      --
    end process;
    -- logger for split-operator array_obj_ref_166_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_166_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_load_0:started:   inputs: " & " valid_1_buffer (guard)= " & Convert_SLV_To_String(valid_1_buffer) & " array_obj_ref_166_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_166_word_address_0));
          --
        end if; 
        if array_obj_ref_166_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_166_load_0:finished:  outputs: " & " array_obj_ref_166_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_166_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_171_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_171_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_load_0:started:   inputs: " & " valid_2_buffer (guard)= " & Convert_SLV_To_String(valid_2_buffer) & " array_obj_ref_171_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_171_word_address_0));
          --
        end if; 
        if array_obj_ref_171_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_171_load_0:finished:  outputs: " & " array_obj_ref_171_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_171_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_166_load_0 array_obj_ref_171_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_166_load_0_req_0,
        array_obj_ref_166_load_0_ack_0,
        array_obj_ref_166_load_0_req_1,
        array_obj_ref_166_load_0_ack_1,
        "array_obj_ref_166_load_0",
        "memory_space_1" ,
        array_obj_ref_166_data_0,
        array_obj_ref_166_word_address_0,
        "array_obj_ref_166_data_0",
        "array_obj_ref_166_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_171_load_0_req_0,
        array_obj_ref_171_load_0_ack_0,
        array_obj_ref_171_load_0_req_1,
        array_obj_ref_171_load_0_ack_1,
        "array_obj_ref_171_load_0",
        "memory_space_1" ,
        array_obj_ref_171_data_0,
        array_obj_ref_171_word_address_0,
        "array_obj_ref_171_data_0",
        "array_obj_ref_171_word_address_0" -- 
      );
      reqL_unguarded(1) <= array_obj_ref_166_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_171_load_0_req_0;
      array_obj_ref_166_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_171_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= array_obj_ref_166_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_171_load_0_req_1;
      array_obj_ref_166_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_171_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= valid_2_buffer(0);
      guard_vector(1)  <= valid_1_buffer(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_166_word_address_0 & array_obj_ref_171_word_address_0;
      array_obj_ref_166_data_0 <= data_out(63 downto 32);
      array_obj_ref_171_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(5 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator array_obj_ref_193_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_193_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_store_0:started:   inputs: " & " valid_w_buffer (guard)= " & Convert_SLV_To_String(valid_w_buffer) & " array_obj_ref_193_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_193_word_address_0) & " array_obj_ref_193_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_193_data_0));
          --
        end if; 
        if array_obj_ref_193_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessReg:DP:array_obj_ref_193_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_193_store_0_req_0,
      array_obj_ref_193_store_0_ack_0,
      array_obj_ref_193_store_0_req_1,
      array_obj_ref_193_store_0_ack_1,
      "array_obj_ref_193_store_0",
      "memory_space_1" ,
      array_obj_ref_193_data_0,
      array_obj_ref_193_word_address_0,
      "array_obj_ref_193_data_0",
      "array_obj_ref_193_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_193_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_193_store_0_req_0;
      array_obj_ref_193_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_193_store_0_req_1;
      array_obj_ref_193_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= valid_w_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_193_word_address_0;
      data_in <= array_obj_ref_193_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(5 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessReg_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity iExecStage is -- 
  generic (tag_length : integer); 
  port ( -- 
    iexec_state : in  std_logic_vector(105 downto 0);
    iexec_rd1_final : in  std_logic_vector(31 downto 0);
    iexec_rd2_final : in  std_logic_vector(31 downto 0);
    next_dcache_state : out  std_logic_vector(138 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity iExecStage;
architecture iExecStage_arch of iExecStage is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 170)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 139)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal iexec_state_buffer :  std_logic_vector(105 downto 0);
  signal iexec_state_update_enable: Boolean;
  signal iexec_rd1_final_buffer :  std_logic_vector(31 downto 0);
  signal iexec_rd1_final_update_enable: Boolean;
  signal iexec_rd2_final_buffer :  std_logic_vector(31 downto 0);
  signal iexec_rd2_final_update_enable: Boolean;
  -- output port buffer signals
  signal next_dcache_state_buffer :  std_logic_vector(138 downto 0);
  signal next_dcache_state_update_enable: Boolean;
  signal iExecStage_CP_456_start: Boolean;
  signal iExecStage_CP_456_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_0 : boolean;
  signal OR_u32_u32_292_inst_req_1 : boolean;
  signal W_is_rs1_neg_404_delayed_1_0_436_inst_ack_0 : boolean;
  signal NOT_u1_u1_434_inst_ack_1 : boolean;
  signal NOT_u1_u1_434_inst_req_1 : boolean;
  signal NOT_u1_u1_434_inst_ack_0 : boolean;
  signal NOT_u1_u1_434_inst_req_0 : boolean;
  signal ADD_u32_u32_253_inst_ack_0 : boolean;
  signal OR_u32_u32_292_inst_ack_0 : boolean;
  signal OR_u32_u32_292_inst_req_0 : boolean;
  signal AND_u32_u32_238_inst_ack_1 : boolean;
  signal W_iexec_rd2_final_418_delayed_1_0_455_inst_req_0 : boolean;
  signal XOR_u32_u32_243_inst_ack_1 : boolean;
  signal type_cast_270_inst_ack_0 : boolean;
  signal XOR_u32_u32_243_inst_req_1 : boolean;
  signal type_cast_270_inst_req_0 : boolean;
  signal XOR_u32_u32_243_inst_ack_0 : boolean;
  signal XOR_u32_u32_243_inst_req_0 : boolean;
  signal type_cast_264_inst_ack_0 : boolean;
  signal type_cast_264_inst_req_0 : boolean;
  signal XOR_u32_u32_248_inst_req_1 : boolean;
  signal AND_u32_u32_238_inst_req_1 : boolean;
  signal AND_u32_u32_238_inst_ack_0 : boolean;
  signal AND_u32_u32_238_inst_req_0 : boolean;
  signal W_iexec_rd1_final_357_delayed_1_0_386_inst_req_0 : boolean;
  signal ADD_u32_u32_253_inst_ack_1 : boolean;
  signal OR_u32_u32_233_inst_ack_1 : boolean;
  signal OR_u32_u32_233_inst_req_1 : boolean;
  signal W_is_rs1_neg_404_delayed_1_0_436_inst_req_1 : boolean;
  signal SUB_u32_u32_258_inst_req_0 : boolean;
  signal type_cast_270_inst_ack_1 : boolean;
  signal ADD_u32_u32_253_inst_req_1 : boolean;
  signal slice_207_inst_req_0 : boolean;
  signal SUB_u32_u32_258_inst_ack_0 : boolean;
  signal W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_0 : boolean;
  signal W_iexec_rd1_final_364_delayed_1_0_398_inst_req_0 : boolean;
  signal W_iexec_rd1_final_357_delayed_1_0_386_inst_req_1 : boolean;
  signal W_iexec_rd2_final_369_delayed_1_0_401_inst_req_0 : boolean;
  signal slice_211_inst_req_1 : boolean;
  signal slice_215_inst_ack_0 : boolean;
  signal slice_215_inst_req_0 : boolean;
  signal W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_1 : boolean;
  signal slice_211_inst_ack_0 : boolean;
  signal slice_211_inst_req_0 : boolean;
  signal type_cast_264_inst_ack_1 : boolean;
  signal W_iexec_rd1_final_364_delayed_1_0_398_inst_req_1 : boolean;
  signal type_cast_264_inst_req_1 : boolean;
  signal W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_1 : boolean;
  signal W_iexec_rd2_final_369_delayed_1_0_401_inst_req_1 : boolean;
  signal W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_0 : boolean;
  signal W_iexec_rd1_final_415_delayed_1_0_452_inst_req_1 : boolean;
  signal W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_1 : boolean;
  signal CONCAT_u64_u139_475_inst_req_0 : boolean;
  signal W_iexec_rd2_final_418_delayed_1_0_455_inst_req_1 : boolean;
  signal W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_1 : boolean;
  signal ADD_u32_u32_253_inst_req_0 : boolean;
  signal XOR_u32_u32_248_inst_ack_1 : boolean;
  signal OR_u32_u32_233_inst_ack_0 : boolean;
  signal type_cast_270_inst_req_1 : boolean;
  signal W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_1 : boolean;
  signal W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_0 : boolean;
  signal OR_u32_u32_233_inst_req_0 : boolean;
  signal AND_u32_u32_228_inst_ack_1 : boolean;
  signal AND_u32_u32_228_inst_req_1 : boolean;
  signal AND_u32_u32_228_inst_ack_0 : boolean;
  signal W_iexec_rd1_final_415_delayed_1_0_452_inst_req_0 : boolean;
  signal W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_0 : boolean;
  signal AND_u32_u32_228_inst_req_0 : boolean;
  signal slice_223_inst_ack_1 : boolean;
  signal slice_223_inst_req_1 : boolean;
  signal slice_223_inst_ack_0 : boolean;
  signal OR_u32_u32_292_inst_ack_1 : boolean;
  signal slice_223_inst_req_0 : boolean;
  signal slice_207_inst_ack_1 : boolean;
  signal SUB_u32_u32_258_inst_ack_1 : boolean;
  signal W_is_rs1_neg_404_delayed_1_0_436_inst_ack_1 : boolean;
  signal slice_219_inst_ack_1 : boolean;
  signal slice_219_inst_req_1 : boolean;
  signal SUB_u32_u32_258_inst_req_1 : boolean;
  signal slice_219_inst_ack_0 : boolean;
  signal slice_219_inst_req_0 : boolean;
  signal XOR_u32_u32_248_inst_ack_0 : boolean;
  signal slice_215_inst_req_1 : boolean;
  signal W_is_rs1_neg_404_delayed_1_0_436_inst_req_0 : boolean;
  signal XOR_u32_u32_248_inst_req_0 : boolean;
  signal slice_215_inst_ack_1 : boolean;
  signal W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_1 : boolean;
  signal W_iexec_rd2_final_358_delayed_1_0_389_inst_req_1 : boolean;
  signal W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_0 : boolean;
  signal W_iexec_rd2_final_358_delayed_1_0_389_inst_req_0 : boolean;
  signal slice_207_inst_req_1 : boolean;
  signal slice_211_inst_ack_1 : boolean;
  signal slice_207_inst_ack_0 : boolean;
  signal CONCAT_u64_u139_475_inst_ack_0 : boolean;
  signal CONCAT_u64_u139_475_inst_req_1 : boolean;
  signal CONCAT_u64_u139_475_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "iExecStage_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 170) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(105 downto 0) <= iexec_state;
  iexec_state_buffer <= in_buffer_data_out(105 downto 0);
  in_buffer_data_in(137 downto 106) <= iexec_rd1_final;
  iexec_rd1_final_buffer <= in_buffer_data_out(137 downto 106);
  in_buffer_data_in(169 downto 138) <= iexec_rd2_final;
  iexec_rd2_final_buffer <= in_buffer_data_out(169 downto 138);
  in_buffer_data_in(tag_length + 169 downto 170) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 169 downto 170);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 1,4 => 7);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 7);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= iexec_state_update_enable & iexec_rd1_final_update_enable & iexec_rd2_final_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  iExecStage_CP_456_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "iExecStage_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 139) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(138 downto 0) <= next_dcache_state_buffer;
  next_dcache_state <= out_buffer_data_out(138 downto 0);
  out_buffer_data_in(tag_length + 138 downto 139) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 138 downto 139);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= iExecStage_CP_456_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  next_dcache_state_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 36) := "next_dcache_state_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_next_dcache_state_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => next_dcache_state_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= iExecStage_CP_456_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= iExecStage_CP_456_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,iExecStage_CP_456_start,"iExecStage cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,iExecStage_CP_456_symbol, "iExecStage cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  iExecStage_CP_456: Block -- control-path 
    signal iExecStage_CP_456_elements: BooleanArray(106 downto 0);
    -- 
  begin -- 
    iExecStage_CP_456_elements(0) <= iExecStage_CP_456_start;
    iExecStage_CP_456_symbol <= iExecStage_CP_456_elements(106);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	22 
    -- CP-element group 1: 	26 
    -- CP-element group 1: 	30 
    -- CP-element group 1: 	34 
    -- CP-element group 1: 	38 
    -- CP-element group 1: 	42 
    -- CP-element group 1: 	46 
    -- CP-element group 1: 	50 
    -- CP-element group 1: 	54 
    -- CP-element group 1: 	58 
    -- CP-element group 1: 	62 
    -- CP-element group 1: 	66 
    -- CP-element group 1: 	70 
    -- CP-element group 1: 	74 
    -- CP-element group 1: 	78 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_208_to_assign_stmt_476/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_CP_456_elements(1) <= iExecStage_CP_456_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	24 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	102 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_476/iexec_state_update_enable_out
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_476/iexec_state_update_enable
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "iExecStage_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(8) & iExecStage_CP_456_elements(12) & iExecStage_CP_456_elements(16) & iExecStage_CP_456_elements(20) & iExecStage_CP_456_elements(24);
      gj_iExecStage_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	28 
    -- CP-element group 3: 	32 
    -- CP-element group 3: 	40 
    -- CP-element group 3: 	44 
    -- CP-element group 3: 	48 
    -- CP-element group 3: 	52 
    -- CP-element group 3: 	56 
    -- CP-element group 3: 	60 
    -- CP-element group 3: 	64 
    -- CP-element group 3: 	68 
    -- CP-element group 3: 	76 
    -- CP-element group 3: 	84 
    -- CP-element group 3: 	88 
    -- CP-element group 3: 	92 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	103 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_208_to_assign_stmt_476/iexec_rd1_final_update_enable_out
      -- CP-element group 3: 	 assign_stmt_208_to_assign_stmt_476/iexec_rd1_final_update_enable
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 29) := "iExecStage_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(28) & iExecStage_CP_456_elements(32) & iExecStage_CP_456_elements(40) & iExecStage_CP_456_elements(44) & iExecStage_CP_456_elements(48) & iExecStage_CP_456_elements(52) & iExecStage_CP_456_elements(56) & iExecStage_CP_456_elements(60) & iExecStage_CP_456_elements(64) & iExecStage_CP_456_elements(68) & iExecStage_CP_456_elements(76) & iExecStage_CP_456_elements(84) & iExecStage_CP_456_elements(88) & iExecStage_CP_456_elements(92);
      gj_iExecStage_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	28 
    -- CP-element group 4: 	32 
    -- CP-element group 4: 	36 
    -- CP-element group 4: 	40 
    -- CP-element group 4: 	44 
    -- CP-element group 4: 	48 
    -- CP-element group 4: 	52 
    -- CP-element group 4: 	56 
    -- CP-element group 4: 	60 
    -- CP-element group 4: 	64 
    -- CP-element group 4: 	72 
    -- CP-element group 4: 	80 
    -- CP-element group 4: 	96 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	104 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_208_to_assign_stmt_476/iexec_rd2_final_update_enable_out
      -- CP-element group 4: 	 assign_stmt_208_to_assign_stmt_476/iexec_rd2_final_update_enable
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 29) := "iExecStage_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(28) & iExecStage_CP_456_elements(32) & iExecStage_CP_456_elements(36) & iExecStage_CP_456_elements(40) & iExecStage_CP_456_elements(44) & iExecStage_CP_456_elements(48) & iExecStage_CP_456_elements(52) & iExecStage_CP_456_elements(56) & iExecStage_CP_456_elements(60) & iExecStage_CP_456_elements(64) & iExecStage_CP_456_elements(72) & iExecStage_CP_456_elements(80) & iExecStage_CP_456_elements(96);
      gj_iExecStage_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	105 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	99 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_208_to_assign_stmt_476/next_dcache_state_update_enable
      -- CP-element group 5: 	 assign_stmt_208_to_assign_stmt_476/next_dcache_state_update_enable_in
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_CP_456_elements(5) <= iExecStage_CP_456_elements(105);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_208_to_assign_stmt_476/slice_207_sample_start_
      -- CP-element group 6: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Sample/rr
      -- CP-element group 6: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Sample/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_207_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(6), ack => slice_207_inst_req_0); -- 
    iExecStage_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "iExecStage_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(8);
      gj_iExecStage_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: 	100 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Update/cr
      -- CP-element group 7: 	 assign_stmt_208_to_assign_stmt_476/slice_207_update_start_
      -- CP-element group 7: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_207_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(7), ack => slice_207_inst_req_1); -- 
    iExecStage_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "iExecStage_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(9) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_208_to_assign_stmt_476/slice_207_sample_completed_
      -- CP-element group 8: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Sample/ra
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_207_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_207_inst_ack_0, ack => iExecStage_CP_456_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	98 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_208_to_assign_stmt_476/slice_207_update_completed_
      -- CP-element group 9: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Update/ca
      -- CP-element group 9: 	 assign_stmt_208_to_assign_stmt_476/slice_207_Update/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_207_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_207_inst_ack_1, ack => iExecStage_CP_456_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Sample/rr
      -- CP-element group 10: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_208_to_assign_stmt_476/slice_211_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_211_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(10), ack => slice_211_inst_req_0); -- 
    iExecStage_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(12);
      gj_iExecStage_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: 	100 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Update/cr
      -- CP-element group 11: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Update/$entry
      -- CP-element group 11: 	 assign_stmt_208_to_assign_stmt_476/slice_211_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_211_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(11), ack => slice_211_inst_req_1); -- 
    iExecStage_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(13) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Sample/ra
      -- CP-element group 12: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_208_to_assign_stmt_476/slice_211_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_211_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_211_inst_ack_0, ack => iExecStage_CP_456_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	98 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Update/$exit
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_476/slice_211_update_completed_
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_476/slice_211_Update/ca
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_211_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_211_inst_ack_1, ack => iExecStage_CP_456_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Sample/rr
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_476/slice_215_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_215_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(14), ack => slice_215_inst_req_0); -- 
    iExecStage_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(16);
      gj_iExecStage_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	100 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Update/$entry
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Update/cr
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_476/slice_215_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_215_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(15), ack => slice_215_inst_req_1); -- 
    iExecStage_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(17) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Sample/ra
      -- CP-element group 16: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_208_to_assign_stmt_476/slice_215_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_215_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_215_inst_ack_0, ack => iExecStage_CP_456_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	98 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Update/$exit
      -- CP-element group 17: 	 assign_stmt_208_to_assign_stmt_476/slice_215_update_completed_
      -- CP-element group 17: 	 assign_stmt_208_to_assign_stmt_476/slice_215_Update/ca
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_215_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_215_inst_ack_1, ack => iExecStage_CP_456_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Sample/rr
      -- CP-element group 18: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Sample/$entry
      -- CP-element group 18: 	 assign_stmt_208_to_assign_stmt_476/slice_219_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_219_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(18), ack => slice_219_inst_req_0); -- 
    iExecStage_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(20);
      gj_iExecStage_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	100 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Update/cr
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Update/$entry
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_476/slice_219_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_219_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(19), ack => slice_219_inst_req_1); -- 
    iExecStage_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(21) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Sample/ra
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Sample/$exit
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_476/slice_219_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_219_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_219_inst_ack_0, ack => iExecStage_CP_456_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	98 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Update/ca
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_476/slice_219_Update/$exit
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_476/slice_219_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_219_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_219_inst_ack_1, ack => iExecStage_CP_456_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	1 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Sample/rr
      -- CP-element group 22: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_208_to_assign_stmt_476/slice_223_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_223_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(22), ack => slice_223_inst_req_0); -- 
    iExecStage_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(24);
      gj_iExecStage_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	100 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Update/cr
      -- CP-element group 23: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Update/$entry
      -- CP-element group 23: 	 assign_stmt_208_to_assign_stmt_476/slice_223_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_223_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(23), ack => slice_223_inst_req_1); -- 
    iExecStage_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(25) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Sample/ra
      -- CP-element group 24: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_208_to_assign_stmt_476/slice_223_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_223_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_223_inst_ack_0, ack => iExecStage_CP_456_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	98 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Update/ca
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_476/slice_223_Update/$exit
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_476/slice_223_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:slice_223_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_223_inst_ack_1, ack => iExecStage_CP_456_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	1 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Sample/rr
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Sample/$entry
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_228_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(26), ack => AND_u32_u32_228_inst_req_0); -- 
    iExecStage_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(28);
      gj_iExecStage_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	100 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Update/cr
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Update/$entry
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_228_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(27), ack => AND_u32_u32_228_inst_req_1); -- 
    iExecStage_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(29) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	3 
    -- CP-element group 28: 	4 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Sample/ra
      -- CP-element group 28: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Sample/$exit
      -- CP-element group 28: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_228_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_228_inst_ack_0, ack => iExecStage_CP_456_elements(28)); -- 
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	98 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Update/ca
      -- CP-element group 29: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_Update/$exit
      -- CP-element group 29: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_228_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_228_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_228_inst_ack_1, ack => iExecStage_CP_456_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	1 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Sample/rr
      -- CP-element group 30: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_233_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(30), ack => OR_u32_u32_233_inst_req_0); -- 
    iExecStage_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(32);
      gj_iExecStage_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	100 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Update/cr
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Update/$entry
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_233_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(31), ack => OR_u32_u32_233_inst_req_1); -- 
    iExecStage_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(33) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	3 
    -- CP-element group 32: 	4 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Sample/ra
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_233_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_233_inst_ack_0, ack => iExecStage_CP_456_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	98 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Update/ca
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_Update/$exit
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_233_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_233_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_233_inst_ack_1, ack => iExecStage_CP_456_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	1 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Sample/rr
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_238_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(34), ack => AND_u32_u32_238_inst_req_0); -- 
    iExecStage_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(36);
      gj_iExecStage_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	100 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Update/cr
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Update/$entry
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_238_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(35), ack => AND_u32_u32_238_inst_req_1); -- 
    iExecStage_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(37) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	4 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Sample/ra
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Sample/$exit
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_238_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_238_inst_ack_0, ack => iExecStage_CP_456_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	98 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Update/ca
      -- CP-element group 37: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_Update/$exit
      -- CP-element group 37: 	 assign_stmt_208_to_assign_stmt_476/AND_u32_u32_238_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:AND_u32_u32_238_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_238_inst_ack_1, ack => iExecStage_CP_456_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	1 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Sample/rr
      -- CP-element group 38: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Sample/$entry
      -- CP-element group 38: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_243_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(38), ack => XOR_u32_u32_243_inst_req_0); -- 
    iExecStage_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(40);
      gj_iExecStage_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: 	100 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Update/cr
      -- CP-element group 39: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Update/$entry
      -- CP-element group 39: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_243_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(39), ack => XOR_u32_u32_243_inst_req_1); -- 
    iExecStage_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(41) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	3 
    -- CP-element group 40: 	4 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Sample/ra
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Sample/$exit
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_243_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_243_inst_ack_0, ack => iExecStage_CP_456_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	98 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Update/ca
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_Update/$exit
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_243_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_243_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_243_inst_ack_1, ack => iExecStage_CP_456_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	1 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_sample_start_
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Sample/$entry
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Sample/rr
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_248_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(42), ack => XOR_u32_u32_248_inst_req_0); -- 
    iExecStage_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(44);
      gj_iExecStage_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Update/cr
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Update/$entry
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_248_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(43), ack => XOR_u32_u32_248_inst_req_1); -- 
    iExecStage_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(45) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: 	4 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_sample_completed_
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Sample/ra
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Sample/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_248_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_248_inst_ack_0, ack => iExecStage_CP_456_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	98 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	43 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_update_completed_
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Update/$exit
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_476/XOR_u32_u32_248_Update/ca
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:XOR_u32_u32_248_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_248_inst_ack_1, ack => iExecStage_CP_456_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	1 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_sample_start_
      -- CP-element group 46: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Sample/rr
      -- CP-element group 46: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Sample/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:ADD_u32_u32_253_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(46), ack => ADD_u32_u32_253_inst_req_0); -- 
    iExecStage_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(48);
      gj_iExecStage_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Update/cr
      -- CP-element group 47: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_update_start_
      -- CP-element group 47: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:ADD_u32_u32_253_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(47), ack => ADD_u32_u32_253_inst_req_1); -- 
    iExecStage_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(49) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	3 
    -- CP-element group 48: 	4 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Sample/ra
      -- CP-element group 48: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Sample/$exit
      -- CP-element group 48: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:ADD_u32_u32_253_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_253_inst_ack_0, ack => iExecStage_CP_456_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	98 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_update_completed_
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Update/ca
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_476/ADD_u32_u32_253_Update/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:ADD_u32_u32_253_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_253_inst_ack_1, ack => iExecStage_CP_456_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	1 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Sample/rr
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_sample_start_
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Sample/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:SUB_u32_u32_258_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(50), ack => SUB_u32_u32_258_inst_req_0); -- 
    iExecStage_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(52);
      gj_iExecStage_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Update/$entry
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_update_start_
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Update/cr
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:SUB_u32_u32_258_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(51), ack => SUB_u32_u32_258_inst_req_1); -- 
    iExecStage_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(53) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	3 
    -- CP-element group 52: 	4 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_sample_completed_
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Sample/ra
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Sample/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:SUB_u32_u32_258_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_258_inst_ack_0, ack => iExecStage_CP_456_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	98 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_update_completed_
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Update/ca
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_476/SUB_u32_u32_258_Update/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:SUB_u32_u32_258_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_258_inst_ack_1, ack => iExecStage_CP_456_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	1 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Sample/rr
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Sample/$entry
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_264_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(54), ack => type_cast_264_inst_req_0); -- 
    iExecStage_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(56);
      gj_iExecStage_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Update/$entry
      -- CP-element group 55: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_update_start_
      -- CP-element group 55: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Update/cr
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_264_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(55), ack => type_cast_264_inst_req_1); -- 
    iExecStage_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(57) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	3 
    -- CP-element group 56: 	4 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Sample/ra
      -- CP-element group 56: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Sample/$exit
      -- CP-element group 56: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_264_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_0, ack => iExecStage_CP_456_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	98 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	55 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Update/$exit
      -- CP-element group 57: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_update_completed_
      -- CP-element group 57: 	 assign_stmt_208_to_assign_stmt_476/type_cast_264_Update/ca
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_264_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_1, ack => iExecStage_CP_456_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	1 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Sample/rr
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Sample/$entry
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_270_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(58), ack => type_cast_270_inst_req_0); -- 
    iExecStage_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(60);
      gj_iExecStage_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	100 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_update_start_
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Update/cr
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_270_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(59), ack => type_cast_270_inst_req_1); -- 
    iExecStage_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(61) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	3 
    -- CP-element group 60: 	4 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Sample/ra
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Sample/$exit
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_270_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_0, ack => iExecStage_CP_456_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	98 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_update_completed_
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Update/ca
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_476/type_cast_270_Update/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:type_cast_270_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_1, ack => iExecStage_CP_456_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	1 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Sample/$entry
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Sample/rr
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_292_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(62), ack => OR_u32_u32_292_inst_req_0); -- 
    iExecStage_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(64);
      gj_iExecStage_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Update/cr
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Update/$entry
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_292_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(63), ack => OR_u32_u32_292_inst_req_1); -- 
    iExecStage_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(65) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	3 
    -- CP-element group 64: 	4 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Sample/ra
      -- CP-element group 64: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Sample/$exit
      -- CP-element group 64: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_292_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_292_inst_ack_0, ack => iExecStage_CP_456_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	98 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Update/$exit
      -- CP-element group 65: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_update_completed_
      -- CP-element group 65: 	 assign_stmt_208_to_assign_stmt_476/OR_u32_u32_292_Update/ca
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:OR_u32_u32_292_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_292_inst_ack_1, ack => iExecStage_CP_456_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	1 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_sample_start_
      -- CP-element group 66: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Sample/req
      -- CP-element group 66: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Sample/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_357_delayed_1_0_386_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(66), ack => W_iexec_rd1_final_357_delayed_1_0_386_inst_req_0); -- 
    iExecStage_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(68);
      gj_iExecStage_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: 	100 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Update/req
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_update_start_
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_357_delayed_1_0_386_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(67), ack => W_iexec_rd1_final_357_delayed_1_0_386_inst_req_1); -- 
    iExecStage_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(69) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	3 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Sample/ack
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_sample_completed_
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Sample/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_0, ack => iExecStage_CP_456_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	98 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Update/ack
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_update_completed_
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_388_Update/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_1, ack => iExecStage_CP_456_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	1 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Sample/$entry
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_sample_start_
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Sample/req
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_358_delayed_1_0_389_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(70), ack => W_iexec_rd2_final_358_delayed_1_0_389_inst_req_0); -- 
    iExecStage_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(72);
      gj_iExecStage_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	100 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_update_start_
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Update/req
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_358_delayed_1_0_389_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(71), ack => W_iexec_rd2_final_358_delayed_1_0_389_inst_req_1); -- 
    iExecStage_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(73) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	4 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Sample/$exit
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_sample_completed_
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Sample/ack
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_0, ack => iExecStage_CP_456_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	98 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_update_completed_
      -- CP-element group 73: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Update/ack
      -- CP-element group 73: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_391_Update/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_1, ack => iExecStage_CP_456_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	1 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Sample/req
      -- CP-element group 74: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Sample/$entry
      -- CP-element group 74: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_364_delayed_1_0_398_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(74), ack => W_iexec_rd1_final_364_delayed_1_0_398_inst_req_0); -- 
    iExecStage_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(76);
      gj_iExecStage_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	100 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_update_start_
      -- CP-element group 75: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Update/req
      -- CP-element group 75: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_364_delayed_1_0_398_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(75), ack => W_iexec_rd1_final_364_delayed_1_0_398_inst_req_1); -- 
    iExecStage_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(77) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	3 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Sample/ack
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Sample/$exit
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_0, ack => iExecStage_CP_456_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	98 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_update_completed_
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Update/ack
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_400_Update/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_1, ack => iExecStage_CP_456_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	1 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_sample_start_
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Sample/req
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Sample/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_369_delayed_1_0_401_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(78), ack => W_iexec_rd2_final_369_delayed_1_0_401_inst_req_0); -- 
    iExecStage_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(80);
      gj_iExecStage_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: 	100 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Update/req
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Update/$entry
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_369_delayed_1_0_401_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(79), ack => W_iexec_rd2_final_369_delayed_1_0_401_inst_req_1); -- 
    iExecStage_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(81) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	4 
    -- CP-element group 80: 	78 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_sample_completed_
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Sample/ack
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Sample/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_0, ack => iExecStage_CP_456_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	98 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	79 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Update/ack
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_Update/$exit
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_403_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_1, ack => iExecStage_CP_456_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Sample/rr
      -- CP-element group 82: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Sample/$entry
      -- CP-element group 82: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_sample_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:NOT_u1_u1_434_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(82), ack => NOT_u1_u1_434_inst_req_0); -- 
    iExecStage_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(84);
      gj_iExecStage_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: 	100 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Update/cr
      -- CP-element group 83: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Update/$entry
      -- CP-element group 83: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:NOT_u1_u1_434_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(83), ack => NOT_u1_u1_434_inst_req_1); -- 
    iExecStage_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(85) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	3 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Sample/$exit
      -- CP-element group 84: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Sample/ra
      -- CP-element group 84: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_sample_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:NOT_u1_u1_434_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_434_inst_ack_0, ack => iExecStage_CP_456_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	98 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Update/ca
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_Update/$exit
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_476/NOT_u1_u1_434_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:NOT_u1_u1_434_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_434_inst_ack_1, ack => iExecStage_CP_456_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Sample/$entry
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_sample_start_
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Sample/req
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_is_rs1_neg_404_delayed_1_0_436_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(86), ack => W_is_rs1_neg_404_delayed_1_0_436_inst_req_0); -- 
    iExecStage_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(88);
      gj_iExecStage_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: 	100 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Update/req
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_update_start_
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_is_rs1_neg_404_delayed_1_0_436_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(87), ack => W_is_rs1_neg_404_delayed_1_0_436_inst_req_1); -- 
    iExecStage_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(89) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	3 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Sample/ack
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_sample_completed_
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Sample/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_is_rs1_neg_404_delayed_1_0_436_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_rs1_neg_404_delayed_1_0_436_inst_ack_0, ack => iExecStage_CP_456_elements(88)); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	98 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_update_completed_
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Update/$exit
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_438_Update/ack
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_is_rs1_neg_404_delayed_1_0_436_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_rs1_neg_404_delayed_1_0_436_inst_ack_1, ack => iExecStage_CP_456_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_sample_start_
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Sample/req
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Sample/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_415_delayed_1_0_452_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(90), ack => W_iexec_rd1_final_415_delayed_1_0_452_inst_req_0); -- 
    iExecStage_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(92);
      gj_iExecStage_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: 	100 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Update/$entry
      -- CP-element group 91: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Update/req
      -- CP-element group 91: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_update_start_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_415_delayed_1_0_452_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(91), ack => W_iexec_rd1_final_415_delayed_1_0_452_inst_req_1); -- 
    iExecStage_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(93) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	3 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_sample_completed_
      -- CP-element group 92: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Sample/ack
      -- CP-element group 92: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Sample/$exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_0, ack => iExecStage_CP_456_elements(92)); -- 
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	98 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Update/$exit
      -- CP-element group 93: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_Update/ack
      -- CP-element group 93: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_454_update_completed_
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_1, ack => iExecStage_CP_456_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_sample_start_
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Sample/$entry
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Sample/req
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_418_delayed_1_0_455_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(94), ack => W_iexec_rd2_final_418_delayed_1_0_455_inst_req_0); -- 
    iExecStage_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(1) & iExecStage_CP_456_elements(96);
      gj_iExecStage_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	100 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_update_start_
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Update/req
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Update/$entry
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_418_delayed_1_0_455_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(95), ack => W_iexec_rd2_final_418_delayed_1_0_455_inst_req_1); -- 
    iExecStage_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(97) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	4 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_sample_completed_
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Sample/$exit
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Sample/ack
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_0, ack => iExecStage_CP_456_elements(96)); -- 
    -- CP-element group 97:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_update_completed_
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Update/$exit
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_476/assign_stmt_457_Update/ack
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_1, ack => iExecStage_CP_456_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: 	13 
    -- CP-element group 98: 	17 
    -- CP-element group 98: 	21 
    -- CP-element group 98: 	25 
    -- CP-element group 98: 	29 
    -- CP-element group 98: 	33 
    -- CP-element group 98: 	37 
    -- CP-element group 98: 	41 
    -- CP-element group 98: 	45 
    -- CP-element group 98: 	49 
    -- CP-element group 98: 	53 
    -- CP-element group 98: 	57 
    -- CP-element group 98: 	61 
    -- CP-element group 98: 	65 
    -- CP-element group 98: 	69 
    -- CP-element group 98: 	73 
    -- CP-element group 98: 	77 
    -- CP-element group 98: 	81 
    -- CP-element group 98: 	85 
    -- CP-element group 98: 	89 
    -- CP-element group 98: 	93 
    -- CP-element group 98: 	97 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_sample_start_
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Sample/$entry
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Sample/rr
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:CONCAT_u64_u139_475_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(98), ack => CONCAT_u64_u139_475_inst_req_0); -- 
    iExecStage_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 23) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1);
      constant place_markings: IntegerArray(0 to 23)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 1);
      constant place_delays: IntegerArray(0 to 23) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 1);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 24); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(9) & iExecStage_CP_456_elements(13) & iExecStage_CP_456_elements(17) & iExecStage_CP_456_elements(21) & iExecStage_CP_456_elements(25) & iExecStage_CP_456_elements(29) & iExecStage_CP_456_elements(33) & iExecStage_CP_456_elements(37) & iExecStage_CP_456_elements(41) & iExecStage_CP_456_elements(45) & iExecStage_CP_456_elements(49) & iExecStage_CP_456_elements(53) & iExecStage_CP_456_elements(57) & iExecStage_CP_456_elements(61) & iExecStage_CP_456_elements(65) & iExecStage_CP_456_elements(69) & iExecStage_CP_456_elements(73) & iExecStage_CP_456_elements(77) & iExecStage_CP_456_elements(81) & iExecStage_CP_456_elements(85) & iExecStage_CP_456_elements(89) & iExecStage_CP_456_elements(93) & iExecStage_CP_456_elements(97) & iExecStage_CP_456_elements(100);
      gj_iExecStage_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 24, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	5 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_update_start_
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Update/$entry
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Update/cr
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:CONCAT_u64_u139_475_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iExecStage_CP_456_elements(99), ack => CONCAT_u64_u139_475_inst_req_1); -- 
    iExecStage_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "iExecStage_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iExecStage_CP_456_elements(5) & iExecStage_CP_456_elements(101);
      gj_iExecStage_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iExecStage_CP_456_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	7 
    -- CP-element group 100: 	11 
    -- CP-element group 100: 	15 
    -- CP-element group 100: 	19 
    -- CP-element group 100: 	23 
    -- CP-element group 100: 	27 
    -- CP-element group 100: 	31 
    -- CP-element group 100: 	35 
    -- CP-element group 100: 	39 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	59 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	67 
    -- CP-element group 100: 	71 
    -- CP-element group 100: 	75 
    -- CP-element group 100: 	79 
    -- CP-element group 100: 	83 
    -- CP-element group 100: 	87 
    -- CP-element group 100: 	91 
    -- CP-element group 100: 	95 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_sample_completed_
      -- CP-element group 100: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Sample/$exit
      -- CP-element group 100: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Sample/ra
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:CONCAT_u64_u139_475_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u139_475_inst_ack_0, ack => iExecStage_CP_456_elements(100)); -- 
    -- CP-element group 101:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	106 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	99 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 assign_stmt_208_to_assign_stmt_476/$exit
      -- CP-element group 101: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_update_completed_
      -- CP-element group 101: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Update/$exit
      -- CP-element group 101: 	 assign_stmt_208_to_assign_stmt_476/CONCAT_u64_u139_475_Update/ca
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:CONCAT_u64_u139_475_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u139_475_inst_ack_1, ack => iExecStage_CP_456_elements(101)); -- 
    -- CP-element group 102:  place  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	2 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 iexec_state_update_enable
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(102) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_CP_456_elements(102) <= iExecStage_CP_456_elements(2);
    -- CP-element group 103:  place  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	3 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 iexec_rd1_final_update_enable
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(103) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_CP_456_elements(103) <= iExecStage_CP_456_elements(3);
    -- CP-element group 104:  place  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	4 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 iexec_rd2_final_update_enable
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(104) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_CP_456_elements(104) <= iExecStage_CP_456_elements(4);
    -- CP-element group 105:  place  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	5 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 next_dcache_state_update_enable
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(105) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 106:  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	101 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 $exit
      -- 
    -- logger for CP element group iExecStage_CP_456_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and iExecStage_CP_456_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:iExecStage:CP:iExecStage_CP_456_elements(106) fired."); 
        -- 
      end if; --
    end process; 
    iExecStage_CP_456_elements(106) <= iExecStage_CP_456_elements(101);
    --  hookup: inputs to control-path 
    iExecStage_CP_456_elements(105) <= next_dcache_state_update_enable;
    -- hookup: output from control-path 
    iexec_state_update_enable <= iExecStage_CP_456_elements(102);
    iexec_rd1_final_update_enable <= iExecStage_CP_456_elements(103);
    iexec_rd2_final_update_enable <= iExecStage_CP_456_elements(104);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u10_u10_370_wire : std_logic_vector(9 downto 0);
    signal ADD_u32_u32_276_276_delayed_1_0_254 : std_logic_vector(31 downto 0);
    signal AND_u1_u1_444_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_449_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_230_230_delayed_1_0_239 : std_logic_vector(31 downto 0);
    signal AND_u32_u32_241_241_delayed_1_0_229 : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u24_463_wire : std_logic_vector(23 downto 0);
    signal CONCAT_u1_u11_473_wire : std_logic_vector(10 downto 0);
    signal CONCAT_u24_u64_467_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_470_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u64_u75_474_wire : std_logic_vector(74 downto 0);
    signal CONCAT_u8_u16_461_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u40_466_wire : std_logic_vector(39 downto 0);
    signal EQ_u32_u1_275_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_297_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_306_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_313_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_320_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_326_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_333_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_341_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_347_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_354_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_361_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_367_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_381_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_442_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_447_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_269_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_409_wire : std_logic_vector(31 downto 0);
    signal MUX_278_wire : std_logic_vector(31 downto 0);
    signal MUX_284_wire : std_logic_vector(31 downto 0);
    signal MUX_291_wire : std_logic_vector(31 downto 0);
    signal MUX_303_wire : std_logic_vector(31 downto 0);
    signal MUX_309_wire : std_logic_vector(31 downto 0);
    signal MUX_316_wire : std_logic_vector(31 downto 0);
    signal MUX_323_wire : std_logic_vector(31 downto 0);
    signal MUX_329_wire : std_logic_vector(31 downto 0);
    signal MUX_336_wire : std_logic_vector(31 downto 0);
    signal MUX_344_wire : std_logic_vector(31 downto 0);
    signal MUX_350_wire : std_logic_vector(31 downto 0);
    signal MUX_357_wire : std_logic_vector(31 downto 0);
    signal MUX_364_wire : std_logic_vector(31 downto 0);
    signal MUX_373_wire : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_399_399_delayed_1_0_435 : std_logic_vector(0 downto 0);
    signal OR_u32_u32_250_250_delayed_1_0_234 : std_logic_vector(31 downto 0);
    signal OR_u32_u32_285_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_301_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_310_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_317_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_330_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_331_331_delayed_1_0_293 : std_logic_vector(31 downto 0);
    signal OR_u32_u32_337_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_338_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_351_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_358_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_374_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_375_wire : std_logic_vector(31 downto 0);
    signal R_ADD_332_wire_constant : std_logic_vector(7 downto 0);
    signal R_BN_446_wire_constant : std_logic_vector(7 downto 0);
    signal R_BZ_441_wire_constant : std_logic_vector(7 downto 0);
    signal R_CALL_366_wire_constant : std_logic_vector(7 downto 0);
    signal R_CMP_360_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_AND_305_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_OR_312_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SLL_346_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SRA_380_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SRL_353_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_XNOR_319_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_XOR_325_wire_constant : std_logic_vector(7 downto 0);
    signal R_SBIR_296_wire_constant : std_logic_vector(7 downto 0);
    signal R_SUB_340_wire_constant : std_logic_vector(7 downto 0);
    signal R_byte_mask_3_bytes_237_wire_constant : std_logic_vector(31 downto 0);
    signal R_minus_1_282_wire_constant : std_logic_vector(31 downto 0);
    signal R_one_1_382_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_32_289_wire_constant : std_logic_vector(31 downto 0);
    signal R_thirty_one_32_408_wire_constant : std_logic_vector(31 downto 0);
    signal R_thirty_two_32_411_wire_constant : std_logic_vector(31 downto 0);
    signal R_zero_1_383_wire_constant : std_logic_vector(0 downto 0);
    signal R_zero_32_276_wire_constant : std_logic_vector(31 downto 0);
    signal R_zero_32_406_wire_constant : std_logic_vector(31 downto 0);
    signal SHL_u32_u32_263_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_286_286_delayed_1_0_259 : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_410_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_413_wire : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_288_wire : std_logic_vector(0 downto 0);
    signal ULT_u32_u1_281_wire : std_logic_vector(0 downto 0);
    signal XOR_u32_u32_259_259_delayed_1_0_244 : std_logic_vector(31 downto 0);
    signal XOR_u32_u32_267_267_delayed_1_0_249 : std_logic_vector(31 downto 0);
    signal bottom_bits_397 : std_logic_vector(31 downto 0);
    signal exec_result_427 : std_logic_vector(31 downto 0);
    signal exec_result_initial_377 : std_logic_vector(31 downto 0);
    signal iexec_rd1_final_357_delayed_1_0_388 : std_logic_vector(31 downto 0);
    signal iexec_rd1_final_364_delayed_1_0_400 : std_logic_vector(31 downto 0);
    signal iexec_rd1_final_415_delayed_1_0_454 : std_logic_vector(31 downto 0);
    signal iexec_rd2_final_358_delayed_1_0_391 : std_logic_vector(31 downto 0);
    signal iexec_rd2_final_369_delayed_1_0_403 : std_logic_vector(31 downto 0);
    signal iexec_rd2_final_418_delayed_1_0_457 : std_logic_vector(31 downto 0);
    signal is_Branch_451 : std_logic_vector(0 downto 0);
    signal is_SRA_385 : std_logic_vector(0 downto 0);
    signal is_rs1_neg_404_delayed_1_0_438 : std_logic_vector(0 downto 0);
    signal is_rs1_neg_431 : std_logic_vector(0 downto 0);
    signal konst_277_wire_constant : std_logic_vector(31 downto 0);
    signal konst_283_wire_constant : std_logic_vector(31 downto 0);
    signal konst_290_wire_constant : std_logic_vector(31 downto 0);
    signal konst_302_wire_constant : std_logic_vector(31 downto 0);
    signal konst_308_wire_constant : std_logic_vector(31 downto 0);
    signal konst_315_wire_constant : std_logic_vector(31 downto 0);
    signal konst_322_wire_constant : std_logic_vector(31 downto 0);
    signal konst_328_wire_constant : std_logic_vector(31 downto 0);
    signal konst_335_wire_constant : std_logic_vector(31 downto 0);
    signal konst_343_wire_constant : std_logic_vector(31 downto 0);
    signal konst_349_wire_constant : std_logic_vector(31 downto 0);
    signal konst_356_wire_constant : std_logic_vector(31 downto 0);
    signal konst_363_wire_constant : std_logic_vector(31 downto 0);
    signal konst_369_wire_constant : std_logic_vector(9 downto 0);
    signal konst_372_wire_constant : std_logic_vector(31 downto 0);
    signal opcode_208 : std_logic_vector(7 downto 0);
    signal program_cnt_224 : std_logic_vector(9 downto 0);
    signal rd_220 : std_logic_vector(7 downto 0);
    signal result_for_SRA_421 : std_logic_vector(31 downto 0);
    signal rs1_imm_212 : std_logic_vector(7 downto 0);
    signal rs2_216 : std_logic_vector(7 downto 0);
    signal top_bits_415 : std_logic_vector(31 downto 0);
    signal type_cast_295_295_delayed_1_0_265 : std_logic_vector(31 downto 0);
    signal type_cast_300_wire : std_logic_vector(31 downto 0);
    signal type_cast_305_305_delayed_1_0_271 : std_logic_vector(31 downto 0);
    signal type_cast_371_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_ADD_332_wire_constant <= "00001001";
    R_BN_446_wire_constant <= "00001111";
    R_BZ_441_wire_constant <= "00001110";
    R_CALL_366_wire_constant <= "00010000";
    R_CMP_360_wire_constant <= "00010010";
    R_L_AND_305_wire_constant <= "00000101";
    R_L_OR_312_wire_constant <= "00000110";
    R_L_SLL_346_wire_constant <= "00001011";
    R_L_SRA_380_wire_constant <= "00001101";
    R_L_SRL_353_wire_constant <= "00001100";
    R_L_XNOR_319_wire_constant <= "00000111";
    R_L_XOR_325_wire_constant <= "00001000";
    R_SBIR_296_wire_constant <= "00000010";
    R_SUB_340_wire_constant <= "00001010";
    R_byte_mask_3_bytes_237_wire_constant <= "11111111111111111111111100000000";
    R_minus_1_282_wire_constant <= "11111111111111111111111111111111";
    R_one_1_382_wire_constant <= "1";
    R_one_32_289_wire_constant <= "00000000000000000000000000000001";
    R_thirty_one_32_408_wire_constant <= "00000000000000000000000000011111";
    R_thirty_two_32_411_wire_constant <= "00000000000000000000000000100000";
    R_zero_1_383_wire_constant <= "0";
    R_zero_32_276_wire_constant <= "00000000000000000000000000000000";
    R_zero_32_406_wire_constant <= "00000000000000000000000000000000";
    konst_277_wire_constant <= "00000000000000000000000000000000";
    konst_283_wire_constant <= "00000000000000000000000000000000";
    konst_290_wire_constant <= "00000000000000000000000000000000";
    konst_302_wire_constant <= "00000000000000000000000000000000";
    konst_308_wire_constant <= "00000000000000000000000000000000";
    konst_315_wire_constant <= "00000000000000000000000000000000";
    konst_322_wire_constant <= "00000000000000000000000000000000";
    konst_328_wire_constant <= "00000000000000000000000000000000";
    konst_335_wire_constant <= "00000000000000000000000000000000";
    konst_343_wire_constant <= "00000000000000000000000000000000";
    konst_349_wire_constant <= "00000000000000000000000000000000";
    konst_356_wire_constant <= "00000000000000000000000000000000";
    konst_363_wire_constant <= "00000000000000000000000000000000";
    konst_369_wire_constant <= "0000000001";
    konst_372_wire_constant <= "00000000000000000000000000000000";
    -- logger for split-operator MUX_278_inst flow-through 
    process(MUX_278_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_278_inst:flowthrough inputs: " & " EQ_u32_u1_275_wire = "& Convert_SLV_To_Hex_String(EQ_u32_u1_275_wire) & " R_zero_32_276_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_32_276_wire_constant) & " konst_277_wire_constant = "& Convert_SLV_To_Hex_String(konst_277_wire_constant) & " outputs:" & " MUX_278_wire= "  & Convert_SLV_To_Hex_String(MUX_278_wire));
      --
    end process; 
    -- flow-through select operator MUX_278_inst
    MUX_278_wire <= R_zero_32_276_wire_constant when (EQ_u32_u1_275_wire(0) /=  '0') else konst_277_wire_constant;
    -- logger for split-operator MUX_284_inst flow-through 
    process(MUX_284_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_284_inst:flowthrough inputs: " & " ULT_u32_u1_281_wire = "& Convert_SLV_To_Hex_String(ULT_u32_u1_281_wire) & " R_minus_1_282_wire_constant = "& Convert_SLV_To_Hex_String(R_minus_1_282_wire_constant) & " konst_283_wire_constant = "& Convert_SLV_To_Hex_String(konst_283_wire_constant) & " outputs:" & " MUX_284_wire= "  & Convert_SLV_To_Hex_String(MUX_284_wire));
      --
    end process; 
    -- flow-through select operator MUX_284_inst
    MUX_284_wire <= R_minus_1_282_wire_constant when (ULT_u32_u1_281_wire(0) /=  '0') else konst_283_wire_constant;
    -- logger for split-operator MUX_291_inst flow-through 
    process(MUX_291_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_291_inst:flowthrough inputs: " & " UGT_u32_u1_288_wire = "& Convert_SLV_To_Hex_String(UGT_u32_u1_288_wire) & " R_one_32_289_wire_constant = "& Convert_SLV_To_Hex_String(R_one_32_289_wire_constant) & " konst_290_wire_constant = "& Convert_SLV_To_Hex_String(konst_290_wire_constant) & " outputs:" & " MUX_291_wire= "  & Convert_SLV_To_Hex_String(MUX_291_wire));
      --
    end process; 
    -- flow-through select operator MUX_291_inst
    MUX_291_wire <= R_one_32_289_wire_constant when (UGT_u32_u1_288_wire(0) /=  '0') else konst_290_wire_constant;
    -- logger for split-operator MUX_303_inst flow-through 
    process(MUX_303_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_303_inst:flowthrough inputs: " & " EQ_u8_u1_297_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_297_wire) & " OR_u32_u32_301_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_301_wire) & " konst_302_wire_constant = "& Convert_SLV_To_Hex_String(konst_302_wire_constant) & " outputs:" & " MUX_303_wire= "  & Convert_SLV_To_Hex_String(MUX_303_wire));
      --
    end process; 
    -- flow-through select operator MUX_303_inst
    MUX_303_wire <= OR_u32_u32_301_wire when (EQ_u8_u1_297_wire(0) /=  '0') else konst_302_wire_constant;
    -- logger for split-operator MUX_309_inst flow-through 
    process(MUX_309_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_309_inst:flowthrough inputs: " & " EQ_u8_u1_306_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_306_wire) & " AND_u32_u32_241_241_delayed_1_0_229 = "& Convert_SLV_To_Hex_String(AND_u32_u32_241_241_delayed_1_0_229) & " konst_308_wire_constant = "& Convert_SLV_To_Hex_String(konst_308_wire_constant) & " outputs:" & " MUX_309_wire= "  & Convert_SLV_To_Hex_String(MUX_309_wire));
      --
    end process; 
    -- flow-through select operator MUX_309_inst
    MUX_309_wire <= AND_u32_u32_241_241_delayed_1_0_229 when (EQ_u8_u1_306_wire(0) /=  '0') else konst_308_wire_constant;
    -- logger for split-operator MUX_316_inst flow-through 
    process(MUX_316_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_316_inst:flowthrough inputs: " & " EQ_u8_u1_313_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_313_wire) & " OR_u32_u32_250_250_delayed_1_0_234 = "& Convert_SLV_To_Hex_String(OR_u32_u32_250_250_delayed_1_0_234) & " konst_315_wire_constant = "& Convert_SLV_To_Hex_String(konst_315_wire_constant) & " outputs:" & " MUX_316_wire= "  & Convert_SLV_To_Hex_String(MUX_316_wire));
      --
    end process; 
    -- flow-through select operator MUX_316_inst
    MUX_316_wire <= OR_u32_u32_250_250_delayed_1_0_234 when (EQ_u8_u1_313_wire(0) /=  '0') else konst_315_wire_constant;
    -- logger for split-operator MUX_323_inst flow-through 
    process(MUX_323_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_323_inst:flowthrough inputs: " & " EQ_u8_u1_320_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_320_wire) & " XOR_u32_u32_259_259_delayed_1_0_244 = "& Convert_SLV_To_Hex_String(XOR_u32_u32_259_259_delayed_1_0_244) & " konst_322_wire_constant = "& Convert_SLV_To_Hex_String(konst_322_wire_constant) & " outputs:" & " MUX_323_wire= "  & Convert_SLV_To_Hex_String(MUX_323_wire));
      --
    end process; 
    -- flow-through select operator MUX_323_inst
    MUX_323_wire <= XOR_u32_u32_259_259_delayed_1_0_244 when (EQ_u8_u1_320_wire(0) /=  '0') else konst_322_wire_constant;
    -- logger for split-operator MUX_329_inst flow-through 
    process(MUX_329_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_329_inst:flowthrough inputs: " & " EQ_u8_u1_326_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_326_wire) & " XOR_u32_u32_267_267_delayed_1_0_249 = "& Convert_SLV_To_Hex_String(XOR_u32_u32_267_267_delayed_1_0_249) & " konst_328_wire_constant = "& Convert_SLV_To_Hex_String(konst_328_wire_constant) & " outputs:" & " MUX_329_wire= "  & Convert_SLV_To_Hex_String(MUX_329_wire));
      --
    end process; 
    -- flow-through select operator MUX_329_inst
    MUX_329_wire <= XOR_u32_u32_267_267_delayed_1_0_249 when (EQ_u8_u1_326_wire(0) /=  '0') else konst_328_wire_constant;
    -- logger for split-operator MUX_336_inst flow-through 
    process(MUX_336_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_336_inst:flowthrough inputs: " & " EQ_u8_u1_333_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_333_wire) & " ADD_u32_u32_276_276_delayed_1_0_254 = "& Convert_SLV_To_Hex_String(ADD_u32_u32_276_276_delayed_1_0_254) & " konst_335_wire_constant = "& Convert_SLV_To_Hex_String(konst_335_wire_constant) & " outputs:" & " MUX_336_wire= "  & Convert_SLV_To_Hex_String(MUX_336_wire));
      --
    end process; 
    -- flow-through select operator MUX_336_inst
    MUX_336_wire <= ADD_u32_u32_276_276_delayed_1_0_254 when (EQ_u8_u1_333_wire(0) /=  '0') else konst_335_wire_constant;
    -- logger for split-operator MUX_344_inst flow-through 
    process(MUX_344_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_344_inst:flowthrough inputs: " & " EQ_u8_u1_341_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_341_wire) & " SUB_u32_u32_286_286_delayed_1_0_259 = "& Convert_SLV_To_Hex_String(SUB_u32_u32_286_286_delayed_1_0_259) & " konst_343_wire_constant = "& Convert_SLV_To_Hex_String(konst_343_wire_constant) & " outputs:" & " MUX_344_wire= "  & Convert_SLV_To_Hex_String(MUX_344_wire));
      --
    end process; 
    -- flow-through select operator MUX_344_inst
    MUX_344_wire <= SUB_u32_u32_286_286_delayed_1_0_259 when (EQ_u8_u1_341_wire(0) /=  '0') else konst_343_wire_constant;
    -- logger for split-operator MUX_350_inst flow-through 
    process(MUX_350_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_350_inst:flowthrough inputs: " & " EQ_u8_u1_347_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_347_wire) & " type_cast_295_295_delayed_1_0_265 = "& Convert_SLV_To_Hex_String(type_cast_295_295_delayed_1_0_265) & " konst_349_wire_constant = "& Convert_SLV_To_Hex_String(konst_349_wire_constant) & " outputs:" & " MUX_350_wire= "  & Convert_SLV_To_Hex_String(MUX_350_wire));
      --
    end process; 
    -- flow-through select operator MUX_350_inst
    MUX_350_wire <= type_cast_295_295_delayed_1_0_265 when (EQ_u8_u1_347_wire(0) /=  '0') else konst_349_wire_constant;
    -- logger for split-operator MUX_357_inst flow-through 
    process(MUX_357_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_357_inst:flowthrough inputs: " & " EQ_u8_u1_354_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_354_wire) & " type_cast_305_305_delayed_1_0_271 = "& Convert_SLV_To_Hex_String(type_cast_305_305_delayed_1_0_271) & " konst_356_wire_constant = "& Convert_SLV_To_Hex_String(konst_356_wire_constant) & " outputs:" & " MUX_357_wire= "  & Convert_SLV_To_Hex_String(MUX_357_wire));
      --
    end process; 
    -- flow-through select operator MUX_357_inst
    MUX_357_wire <= type_cast_305_305_delayed_1_0_271 when (EQ_u8_u1_354_wire(0) /=  '0') else konst_356_wire_constant;
    -- logger for split-operator MUX_364_inst flow-through 
    process(MUX_364_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_364_inst:flowthrough inputs: " & " EQ_u8_u1_361_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_361_wire) & " OR_u32_u32_331_331_delayed_1_0_293 = "& Convert_SLV_To_Hex_String(OR_u32_u32_331_331_delayed_1_0_293) & " konst_363_wire_constant = "& Convert_SLV_To_Hex_String(konst_363_wire_constant) & " outputs:" & " MUX_364_wire= "  & Convert_SLV_To_Hex_String(MUX_364_wire));
      --
    end process; 
    -- flow-through select operator MUX_364_inst
    MUX_364_wire <= OR_u32_u32_331_331_delayed_1_0_293 when (EQ_u8_u1_361_wire(0) /=  '0') else konst_363_wire_constant;
    -- logger for split-operator MUX_373_inst flow-through 
    process(MUX_373_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_373_inst:flowthrough inputs: " & " EQ_u8_u1_367_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_367_wire) & " type_cast_371_wire = "& Convert_SLV_To_Hex_String(type_cast_371_wire) & " konst_372_wire_constant = "& Convert_SLV_To_Hex_String(konst_372_wire_constant) & " outputs:" & " MUX_373_wire= "  & Convert_SLV_To_Hex_String(MUX_373_wire));
      --
    end process; 
    -- flow-through select operator MUX_373_inst
    MUX_373_wire <= type_cast_371_wire when (EQ_u8_u1_367_wire(0) /=  '0') else konst_372_wire_constant;
    -- logger for split-operator MUX_384_inst flow-through 
    process(is_SRA_385) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_384_inst:flowthrough inputs: " & " EQ_u8_u1_381_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_381_wire) & " R_one_1_382_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_382_wire_constant) & " R_zero_1_383_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_1_383_wire_constant) & " outputs:" & " is_SRA_385= "  & Convert_SLV_To_Hex_String(is_SRA_385));
      --
    end process; 
    -- flow-through select operator MUX_384_inst
    is_SRA_385 <= R_one_1_382_wire_constant when (EQ_u8_u1_381_wire(0) /=  '0') else R_zero_1_383_wire_constant;
    -- logger for split-operator MUX_426_inst flow-through 
    process(exec_result_427) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:MUX_426_inst:flowthrough inputs: " & " is_SRA_385 = "& Convert_SLV_To_Hex_String(is_SRA_385) & " result_for_SRA_421 = "& Convert_SLV_To_Hex_String(result_for_SRA_421) & " exec_result_initial_377 = "& Convert_SLV_To_Hex_String(exec_result_initial_377) & " outputs:" & " exec_result_427= "  & Convert_SLV_To_Hex_String(exec_result_427));
      --
    end process; 
    -- flow-through select operator MUX_426_inst
    exec_result_427 <= result_for_SRA_421 when (is_SRA_385(0) /=  '0') else exec_result_initial_377;
    -- logger for split-operator slice_207_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_207_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_207_inst:started:   inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer));
          --
        end if; 
        if slice_207_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_207_inst:finished:  outputs: " & " opcode_208= "  & Convert_SLV_To_Hex_String(opcode_208));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_207_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_207_inst_req_0;
      slice_207_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_207_inst_req_1;
      slice_207_inst_ack_1<= update_ack(0);
      slice_207_inst: SliceSplitProtocol generic map(name => "slice_207_inst", in_data_width => 106, high_index => 105, low_index => 98, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => iexec_state_buffer, dout => opcode_208, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_211_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_211_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_211_inst:started:   inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer));
          --
        end if; 
        if slice_211_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_211_inst:finished:  outputs: " & " rs1_imm_212= "  & Convert_SLV_To_Hex_String(rs1_imm_212));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_211_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_211_inst_req_0;
      slice_211_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_211_inst_req_1;
      slice_211_inst_ack_1<= update_ack(0);
      slice_211_inst: SliceSplitProtocol generic map(name => "slice_211_inst", in_data_width => 106, high_index => 97, low_index => 90, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => iexec_state_buffer, dout => rs1_imm_212, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_215_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_215_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_215_inst:started:   inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer));
          --
        end if; 
        if slice_215_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_215_inst:finished:  outputs: " & " rs2_216= "  & Convert_SLV_To_Hex_String(rs2_216));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_215_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_215_inst_req_0;
      slice_215_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_215_inst_req_1;
      slice_215_inst_ack_1<= update_ack(0);
      slice_215_inst: SliceSplitProtocol generic map(name => "slice_215_inst", in_data_width => 106, high_index => 89, low_index => 82, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => iexec_state_buffer, dout => rs2_216, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_219_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_219_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_219_inst:started:   inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer));
          --
        end if; 
        if slice_219_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_219_inst:finished:  outputs: " & " rd_220= "  & Convert_SLV_To_Hex_String(rd_220));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_219_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_219_inst_req_0;
      slice_219_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_219_inst_req_1;
      slice_219_inst_ack_1<= update_ack(0);
      slice_219_inst: SliceSplitProtocol generic map(name => "slice_219_inst", in_data_width => 106, high_index => 81, low_index => 74, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => iexec_state_buffer, dout => rd_220, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_223_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_223_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_223_inst:started:   inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer));
          --
        end if; 
        if slice_223_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_223_inst:finished:  outputs: " & " program_cnt_224= "  & Convert_SLV_To_Hex_String(program_cnt_224));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_223_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_223_inst_req_0;
      slice_223_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_223_inst_req_1;
      slice_223_inst_ack_1<= update_ack(0);
      slice_223_inst: SliceSplitProtocol generic map(name => "slice_223_inst", in_data_width => 106, high_index => 9, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => iexec_state_buffer, dout => program_cnt_224, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_430_inst flow-through 
    process(is_rs1_neg_431) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:slice_430_inst:flowthrough inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " outputs:" & " is_rs1_neg_431= "  & Convert_SLV_To_Hex_String(is_rs1_neg_431));
      --
    end process; 
    -- flow-through slice operator slice_430_inst
    is_rs1_neg_431 <= iexec_rd1_final_buffer(31 downto 31);
    -- logger for split-operator W_iexec_rd1_final_357_delayed_1_0_386_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd1_final_357_delayed_1_0_386_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer));
          --
        end if; 
        if W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd1_final_357_delayed_1_0_386_inst:finished:  outputs: " & " iexec_rd1_final_357_delayed_1_0_388= "  & Convert_SLV_To_Hex_String(iexec_rd1_final_357_delayed_1_0_388));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iexec_rd1_final_357_delayed_1_0_386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iexec_rd1_final_357_delayed_1_0_386_inst_req_0;
      W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_0<= wack(0);
      rreq(0) <= W_iexec_rd1_final_357_delayed_1_0_386_inst_req_1;
      W_iexec_rd1_final_357_delayed_1_0_386_inst_ack_1<= rack(0);
      W_iexec_rd1_final_357_delayed_1_0_386_inst : InterlockBuffer generic map ( -- 
        name => "W_iexec_rd1_final_357_delayed_1_0_386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iexec_rd1_final_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iexec_rd1_final_357_delayed_1_0_388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iexec_rd1_final_364_delayed_1_0_398_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd1_final_364_delayed_1_0_398_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer));
          --
        end if; 
        if W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd1_final_364_delayed_1_0_398_inst:finished:  outputs: " & " iexec_rd1_final_364_delayed_1_0_400= "  & Convert_SLV_To_Hex_String(iexec_rd1_final_364_delayed_1_0_400));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iexec_rd1_final_364_delayed_1_0_398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iexec_rd1_final_364_delayed_1_0_398_inst_req_0;
      W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_0<= wack(0);
      rreq(0) <= W_iexec_rd1_final_364_delayed_1_0_398_inst_req_1;
      W_iexec_rd1_final_364_delayed_1_0_398_inst_ack_1<= rack(0);
      W_iexec_rd1_final_364_delayed_1_0_398_inst : InterlockBuffer generic map ( -- 
        name => "W_iexec_rd1_final_364_delayed_1_0_398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iexec_rd1_final_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iexec_rd1_final_364_delayed_1_0_400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iexec_rd1_final_415_delayed_1_0_452_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd1_final_415_delayed_1_0_452_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer));
          --
        end if; 
        if W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd1_final_415_delayed_1_0_452_inst:finished:  outputs: " & " iexec_rd1_final_415_delayed_1_0_454= "  & Convert_SLV_To_Hex_String(iexec_rd1_final_415_delayed_1_0_454));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iexec_rd1_final_415_delayed_1_0_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iexec_rd1_final_415_delayed_1_0_452_inst_req_0;
      W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_0<= wack(0);
      rreq(0) <= W_iexec_rd1_final_415_delayed_1_0_452_inst_req_1;
      W_iexec_rd1_final_415_delayed_1_0_452_inst_ack_1<= rack(0);
      W_iexec_rd1_final_415_delayed_1_0_452_inst : InterlockBuffer generic map ( -- 
        name => "W_iexec_rd1_final_415_delayed_1_0_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iexec_rd1_final_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iexec_rd1_final_415_delayed_1_0_454,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iexec_rd2_final_358_delayed_1_0_389_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd2_final_358_delayed_1_0_389_inst:started:   inputs: " & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd2_final_358_delayed_1_0_389_inst:finished:  outputs: " & " iexec_rd2_final_358_delayed_1_0_391= "  & Convert_SLV_To_Hex_String(iexec_rd2_final_358_delayed_1_0_391));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iexec_rd2_final_358_delayed_1_0_389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iexec_rd2_final_358_delayed_1_0_389_inst_req_0;
      W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_0<= wack(0);
      rreq(0) <= W_iexec_rd2_final_358_delayed_1_0_389_inst_req_1;
      W_iexec_rd2_final_358_delayed_1_0_389_inst_ack_1<= rack(0);
      W_iexec_rd2_final_358_delayed_1_0_389_inst : InterlockBuffer generic map ( -- 
        name => "W_iexec_rd2_final_358_delayed_1_0_389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iexec_rd2_final_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iexec_rd2_final_358_delayed_1_0_391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iexec_rd2_final_369_delayed_1_0_401_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd2_final_369_delayed_1_0_401_inst:started:   inputs: " & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd2_final_369_delayed_1_0_401_inst:finished:  outputs: " & " iexec_rd2_final_369_delayed_1_0_403= "  & Convert_SLV_To_Hex_String(iexec_rd2_final_369_delayed_1_0_403));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iexec_rd2_final_369_delayed_1_0_401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iexec_rd2_final_369_delayed_1_0_401_inst_req_0;
      W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_0<= wack(0);
      rreq(0) <= W_iexec_rd2_final_369_delayed_1_0_401_inst_req_1;
      W_iexec_rd2_final_369_delayed_1_0_401_inst_ack_1<= rack(0);
      W_iexec_rd2_final_369_delayed_1_0_401_inst : InterlockBuffer generic map ( -- 
        name => "W_iexec_rd2_final_369_delayed_1_0_401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iexec_rd2_final_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iexec_rd2_final_369_delayed_1_0_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iexec_rd2_final_418_delayed_1_0_455_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd2_final_418_delayed_1_0_455_inst:started:   inputs: " & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_iexec_rd2_final_418_delayed_1_0_455_inst:finished:  outputs: " & " iexec_rd2_final_418_delayed_1_0_457= "  & Convert_SLV_To_Hex_String(iexec_rd2_final_418_delayed_1_0_457));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iexec_rd2_final_418_delayed_1_0_455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iexec_rd2_final_418_delayed_1_0_455_inst_req_0;
      W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_0<= wack(0);
      rreq(0) <= W_iexec_rd2_final_418_delayed_1_0_455_inst_req_1;
      W_iexec_rd2_final_418_delayed_1_0_455_inst_ack_1<= rack(0);
      W_iexec_rd2_final_418_delayed_1_0_455_inst : InterlockBuffer generic map ( -- 
        name => "W_iexec_rd2_final_418_delayed_1_0_455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iexec_rd2_final_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iexec_rd2_final_418_delayed_1_0_457,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_is_rs1_neg_404_delayed_1_0_436_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_is_rs1_neg_404_delayed_1_0_436_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_is_rs1_neg_404_delayed_1_0_436_inst:started:   inputs: " & " is_rs1_neg_431 = "& Convert_SLV_To_Hex_String(is_rs1_neg_431));
          --
        end if; 
        if W_is_rs1_neg_404_delayed_1_0_436_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:W_is_rs1_neg_404_delayed_1_0_436_inst:finished:  outputs: " & " is_rs1_neg_404_delayed_1_0_438= "  & Convert_SLV_To_Hex_String(is_rs1_neg_404_delayed_1_0_438));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_is_rs1_neg_404_delayed_1_0_436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_is_rs1_neg_404_delayed_1_0_436_inst_req_0;
      W_is_rs1_neg_404_delayed_1_0_436_inst_ack_0<= wack(0);
      rreq(0) <= W_is_rs1_neg_404_delayed_1_0_436_inst_req_1;
      W_is_rs1_neg_404_delayed_1_0_436_inst_ack_1<= rack(0);
      W_is_rs1_neg_404_delayed_1_0_436_inst : InterlockBuffer generic map ( -- 
        name => "W_is_rs1_neg_404_delayed_1_0_436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => is_rs1_neg_431,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => is_rs1_neg_404_delayed_1_0_438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_264_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_264_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:type_cast_264_inst:started:   inputs: " & " SHL_u32_u32_263_wire = "& Convert_SLV_To_Hex_String(SHL_u32_u32_263_wire));
          --
        end if; 
        if type_cast_264_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:type_cast_264_inst:finished:  outputs: " & " type_cast_295_295_delayed_1_0_265= "  & Convert_SLV_To_Hex_String(type_cast_295_295_delayed_1_0_265));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_264_inst_req_0;
      type_cast_264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_264_inst_req_1;
      type_cast_264_inst_ack_1<= rack(0);
      type_cast_264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SHL_u32_u32_263_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_295_295_delayed_1_0_265,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_270_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_270_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:type_cast_270_inst:started:   inputs: " & " LSHR_u32_u32_269_wire = "& Convert_SLV_To_Hex_String(LSHR_u32_u32_269_wire));
          --
        end if; 
        if type_cast_270_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:type_cast_270_inst:finished:  outputs: " & " type_cast_305_305_delayed_1_0_271= "  & Convert_SLV_To_Hex_String(type_cast_305_305_delayed_1_0_271));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_270_inst_req_0;
      type_cast_270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_270_inst_req_1;
      type_cast_270_inst_ack_1<= rack(0);
      type_cast_270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => LSHR_u32_u32_269_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_305_305_delayed_1_0_271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_300_inst flow-through 
    process(type_cast_300_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:type_cast_300_inst:flowthrough inputs: " & " rs1_imm_212 = "& Convert_SLV_To_Hex_String(rs1_imm_212) & " outputs:" & " type_cast_300_wire= "  & Convert_SLV_To_Hex_String(type_cast_300_wire));
      --
    end process; 
    -- interlock type_cast_300_inst
    process(rs1_imm_212) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := rs1_imm_212(7 downto 0);
      type_cast_300_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_371_inst flow-through 
    process(type_cast_371_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:type_cast_371_inst:flowthrough inputs: " & " ADD_u10_u10_370_wire = "& Convert_SLV_To_Hex_String(ADD_u10_u10_370_wire) & " outputs:" & " type_cast_371_wire= "  & Convert_SLV_To_Hex_String(type_cast_371_wire));
      --
    end process; 
    -- interlock type_cast_371_inst
    process(ADD_u10_u10_370_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 9 downto 0) := ADD_u10_u10_370_wire(9 downto 0);
      type_cast_371_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ADD_u10_u10_370_inst flow-through 
    process(ADD_u10_u10_370_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:ADD_u10_u10_370_inst:flowthrough inputs: " & " program_cnt_224 = "& Convert_SLV_To_Hex_String(program_cnt_224) & " konst_369_wire_constant = "& Convert_SLV_To_Hex_String(konst_369_wire_constant) & " outputs:" & " ADD_u10_u10_370_wire= "  & Convert_SLV_To_Hex_String(ADD_u10_u10_370_wire));
      --
    end process; 
    -- binary operator ADD_u10_u10_370_inst
    process(program_cnt_224) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApIntAdd_proc(program_cnt_224, konst_369_wire_constant, tmp_var);
      ADD_u10_u10_370_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_253_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u32_u32_253_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:ADD_u32_u32_253_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if ADD_u32_u32_253_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:ADD_u32_u32_253_inst:finished:  outputs: " & " ADD_u32_u32_276_276_delayed_1_0_254= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_276_276_delayed_1_0_254));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : ADD_u32_u32_253_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iexec_rd1_final_buffer & iexec_rd2_final_buffer;
      ADD_u32_u32_276_276_delayed_1_0_254 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_253_inst_req_0;
      ADD_u32_u32_253_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_253_inst_req_1;
      ADD_u32_u32_253_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator AND_u1_u1_444_inst flow-through 
    process(AND_u1_u1_444_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:AND_u1_u1_444_inst:flowthrough inputs: " & " EQ_u8_u1_442_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_442_wire) & " NOT_u1_u1_399_399_delayed_1_0_435 = "& Convert_SLV_To_Hex_String(NOT_u1_u1_399_399_delayed_1_0_435) & " outputs:" & " AND_u1_u1_444_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_444_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_444_inst
    process(EQ_u8_u1_442_wire, NOT_u1_u1_399_399_delayed_1_0_435) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u8_u1_442_wire, NOT_u1_u1_399_399_delayed_1_0_435, tmp_var);
      AND_u1_u1_444_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_449_inst flow-through 
    process(AND_u1_u1_449_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:AND_u1_u1_449_inst:flowthrough inputs: " & " EQ_u8_u1_447_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_447_wire) & " is_rs1_neg_404_delayed_1_0_438 = "& Convert_SLV_To_Hex_String(is_rs1_neg_404_delayed_1_0_438) & " outputs:" & " AND_u1_u1_449_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_449_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_449_inst
    process(EQ_u8_u1_447_wire, is_rs1_neg_404_delayed_1_0_438) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u8_u1_447_wire, is_rs1_neg_404_delayed_1_0_438, tmp_var);
      AND_u1_u1_449_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_228_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if AND_u32_u32_228_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:AND_u32_u32_228_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if AND_u32_u32_228_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:AND_u32_u32_228_inst:finished:  outputs: " & " AND_u32_u32_241_241_delayed_1_0_229= "  & Convert_SLV_To_Hex_String(AND_u32_u32_241_241_delayed_1_0_229));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (4) : AND_u32_u32_228_inst 
    ApIntAnd_group_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iexec_rd1_final_buffer & iexec_rd2_final_buffer;
      AND_u32_u32_241_241_delayed_1_0_229 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_228_inst_req_0;
      AND_u32_u32_228_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_228_inst_req_1;
      AND_u32_u32_228_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- logger for split-operator AND_u32_u32_238_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if AND_u32_u32_238_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:AND_u32_u32_238_inst:started:   inputs: " & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer) & " R_byte_mask_3_bytes_237_wire_constant = "& Convert_SLV_To_Hex_String(R_byte_mask_3_bytes_237_wire_constant));
          --
        end if; 
        if AND_u32_u32_238_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:AND_u32_u32_238_inst:finished:  outputs: " & " AND_u32_u32_230_230_delayed_1_0_239= "  & Convert_SLV_To_Hex_String(AND_u32_u32_230_230_delayed_1_0_239));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (5) : AND_u32_u32_238_inst 
    ApIntAnd_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iexec_rd2_final_buffer;
      AND_u32_u32_230_230_delayed_1_0_239 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_238_inst_req_0;
      AND_u32_u32_238_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_238_inst_req_1;
      AND_u32_u32_238_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_5_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111100000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- logger for split-operator CONCAT_u16_u24_463_inst flow-through 
    process(CONCAT_u16_u24_463_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u16_u24_463_inst:flowthrough inputs: " & " CONCAT_u8_u16_461_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_461_wire) & " rs2_216 = "& Convert_SLV_To_Hex_String(rs2_216) & " outputs:" & " CONCAT_u16_u24_463_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u24_463_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u24_463_inst
    process(CONCAT_u8_u16_461_wire, rs2_216) -- 
      variable tmp_var : std_logic_vector(23 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_461_wire, rs2_216, tmp_var);
      CONCAT_u16_u24_463_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u11_473_inst flow-through 
    process(CONCAT_u1_u11_473_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u1_u11_473_inst:flowthrough inputs: " & " is_Branch_451 = "& Convert_SLV_To_Hex_String(is_Branch_451) & " program_cnt_224 = "& Convert_SLV_To_Hex_String(program_cnt_224) & " outputs:" & " CONCAT_u1_u11_473_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u11_473_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u11_473_inst
    process(is_Branch_451, program_cnt_224) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      ApConcat_proc(is_Branch_451, program_cnt_224, tmp_var);
      CONCAT_u1_u11_473_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u24_u64_467_inst flow-through 
    process(CONCAT_u24_u64_467_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u24_u64_467_inst:flowthrough inputs: " & " CONCAT_u16_u24_463_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u24_463_wire) & " CONCAT_u8_u40_466_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u40_466_wire) & " outputs:" & " CONCAT_u24_u64_467_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u24_u64_467_wire));
      --
    end process; 
    -- binary operator CONCAT_u24_u64_467_inst
    process(CONCAT_u16_u24_463_wire, CONCAT_u8_u40_466_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u24_463_wire, CONCAT_u8_u40_466_wire, tmp_var);
      CONCAT_u24_u64_467_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_470_inst flow-through 
    process(CONCAT_u32_u64_470_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u32_u64_470_inst:flowthrough inputs: " & " iexec_rd2_final_418_delayed_1_0_457 = "& Convert_SLV_To_Hex_String(iexec_rd2_final_418_delayed_1_0_457) & " exec_result_427 = "& Convert_SLV_To_Hex_String(exec_result_427) & " outputs:" & " CONCAT_u32_u64_470_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_470_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_470_inst
    process(iexec_rd2_final_418_delayed_1_0_457, exec_result_427) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(iexec_rd2_final_418_delayed_1_0_457, exec_result_427, tmp_var);
      CONCAT_u32_u64_470_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u64_u139_475_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u64_u139_475_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u64_u139_475_inst:started:   inputs: " & " CONCAT_u24_u64_467_wire = "& Convert_SLV_To_Hex_String(CONCAT_u24_u64_467_wire) & " CONCAT_u64_u75_474_wire = "& Convert_SLV_To_Hex_String(CONCAT_u64_u75_474_wire));
          --
        end if; 
        if CONCAT_u64_u139_475_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u64_u139_475_inst:finished:  outputs: " & " next_dcache_state_buffer= "  & Convert_SLV_To_Hex_String(next_dcache_state_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (10) : CONCAT_u64_u139_475_inst 
    ApConcat_group_10: Block -- 
      signal data_in: std_logic_vector(138 downto 0);
      signal data_out: std_logic_vector(138 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u24_u64_467_wire & CONCAT_u64_u75_474_wire;
      next_dcache_state_buffer <= data_out(138 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u64_u139_475_inst_req_0;
      CONCAT_u64_u139_475_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u64_u139_475_inst_req_1;
      CONCAT_u64_u139_475_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_10_gI: SplitGuardInterface generic map(name => "ApConcat_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 75, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 139,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- logger for split-operator CONCAT_u64_u75_474_inst flow-through 
    process(CONCAT_u64_u75_474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u64_u75_474_inst:flowthrough inputs: " & " CONCAT_u32_u64_470_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_470_wire) & " CONCAT_u1_u11_473_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u11_473_wire) & " outputs:" & " CONCAT_u64_u75_474_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u64_u75_474_wire));
      --
    end process; 
    -- binary operator CONCAT_u64_u75_474_inst
    process(CONCAT_u32_u64_470_wire, CONCAT_u1_u11_473_wire) -- 
      variable tmp_var : std_logic_vector(74 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_470_wire, CONCAT_u1_u11_473_wire, tmp_var);
      CONCAT_u64_u75_474_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u8_u16_461_inst flow-through 
    process(CONCAT_u8_u16_461_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u8_u16_461_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " rs1_imm_212 = "& Convert_SLV_To_Hex_String(rs1_imm_212) & " outputs:" & " CONCAT_u8_u16_461_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_461_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_461_inst
    process(opcode_208, rs1_imm_212) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(opcode_208, rs1_imm_212, tmp_var);
      CONCAT_u8_u16_461_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u8_u40_466_inst flow-through 
    process(CONCAT_u8_u40_466_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:CONCAT_u8_u40_466_inst:flowthrough inputs: " & " rd_220 = "& Convert_SLV_To_Hex_String(rd_220) & " iexec_rd1_final_415_delayed_1_0_454 = "& Convert_SLV_To_Hex_String(iexec_rd1_final_415_delayed_1_0_454) & " outputs:" & " CONCAT_u8_u40_466_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u40_466_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u40_466_inst
    process(rd_220, iexec_rd1_final_415_delayed_1_0_454) -- 
      variable tmp_var : std_logic_vector(39 downto 0); -- 
    begin -- 
      ApConcat_proc(rd_220, iexec_rd1_final_415_delayed_1_0_454, tmp_var);
      CONCAT_u8_u40_466_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_275_inst flow-through 
    process(EQ_u32_u1_275_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u32_u1_275_inst:flowthrough inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer) & " outputs:" & " EQ_u32_u1_275_wire= "  & Convert_SLV_To_Hex_String(EQ_u32_u1_275_wire));
      --
    end process; 
    -- binary operator EQ_u32_u1_275_inst
    process(iexec_rd1_final_buffer, iexec_rd2_final_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iexec_rd1_final_buffer, iexec_rd2_final_buffer, tmp_var);
      EQ_u32_u1_275_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_297_inst flow-through 
    process(EQ_u8_u1_297_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_297_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_SBIR_296_wire_constant = "& Convert_SLV_To_Hex_String(R_SBIR_296_wire_constant) & " outputs:" & " EQ_u8_u1_297_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_297_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_297_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_SBIR_296_wire_constant, tmp_var);
      EQ_u8_u1_297_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_306_inst flow-through 
    process(EQ_u8_u1_306_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_306_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_L_AND_305_wire_constant = "& Convert_SLV_To_Hex_String(R_L_AND_305_wire_constant) & " outputs:" & " EQ_u8_u1_306_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_306_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_306_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_L_AND_305_wire_constant, tmp_var);
      EQ_u8_u1_306_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_313_inst flow-through 
    process(EQ_u8_u1_313_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_313_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_L_OR_312_wire_constant = "& Convert_SLV_To_Hex_String(R_L_OR_312_wire_constant) & " outputs:" & " EQ_u8_u1_313_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_313_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_313_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_L_OR_312_wire_constant, tmp_var);
      EQ_u8_u1_313_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_320_inst flow-through 
    process(EQ_u8_u1_320_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_320_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_L_XNOR_319_wire_constant = "& Convert_SLV_To_Hex_String(R_L_XNOR_319_wire_constant) & " outputs:" & " EQ_u8_u1_320_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_320_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_320_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_L_XNOR_319_wire_constant, tmp_var);
      EQ_u8_u1_320_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_326_inst flow-through 
    process(EQ_u8_u1_326_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_326_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_L_XOR_325_wire_constant = "& Convert_SLV_To_Hex_String(R_L_XOR_325_wire_constant) & " outputs:" & " EQ_u8_u1_326_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_326_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_326_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_L_XOR_325_wire_constant, tmp_var);
      EQ_u8_u1_326_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_333_inst flow-through 
    process(EQ_u8_u1_333_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_333_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_ADD_332_wire_constant = "& Convert_SLV_To_Hex_String(R_ADD_332_wire_constant) & " outputs:" & " EQ_u8_u1_333_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_333_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_333_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_ADD_332_wire_constant, tmp_var);
      EQ_u8_u1_333_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_341_inst flow-through 
    process(EQ_u8_u1_341_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_341_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_SUB_340_wire_constant = "& Convert_SLV_To_Hex_String(R_SUB_340_wire_constant) & " outputs:" & " EQ_u8_u1_341_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_341_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_341_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_SUB_340_wire_constant, tmp_var);
      EQ_u8_u1_341_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_347_inst flow-through 
    process(EQ_u8_u1_347_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_347_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_L_SLL_346_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SLL_346_wire_constant) & " outputs:" & " EQ_u8_u1_347_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_347_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_347_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_L_SLL_346_wire_constant, tmp_var);
      EQ_u8_u1_347_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_354_inst flow-through 
    process(EQ_u8_u1_354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_354_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_L_SRL_353_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SRL_353_wire_constant) & " outputs:" & " EQ_u8_u1_354_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_354_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_354_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_L_SRL_353_wire_constant, tmp_var);
      EQ_u8_u1_354_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_361_inst flow-through 
    process(EQ_u8_u1_361_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_361_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_CMP_360_wire_constant = "& Convert_SLV_To_Hex_String(R_CMP_360_wire_constant) & " outputs:" & " EQ_u8_u1_361_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_361_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_361_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_CMP_360_wire_constant, tmp_var);
      EQ_u8_u1_361_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_367_inst flow-through 
    process(EQ_u8_u1_367_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_367_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_CALL_366_wire_constant = "& Convert_SLV_To_Hex_String(R_CALL_366_wire_constant) & " outputs:" & " EQ_u8_u1_367_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_367_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_367_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_CALL_366_wire_constant, tmp_var);
      EQ_u8_u1_367_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_381_inst flow-through 
    process(EQ_u8_u1_381_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_381_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_L_SRA_380_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SRA_380_wire_constant) & " outputs:" & " EQ_u8_u1_381_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_381_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_381_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_L_SRA_380_wire_constant, tmp_var);
      EQ_u8_u1_381_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_442_inst flow-through 
    process(EQ_u8_u1_442_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_442_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_BZ_441_wire_constant = "& Convert_SLV_To_Hex_String(R_BZ_441_wire_constant) & " outputs:" & " EQ_u8_u1_442_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_442_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_442_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_BZ_441_wire_constant, tmp_var);
      EQ_u8_u1_442_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_447_inst flow-through 
    process(EQ_u8_u1_447_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:EQ_u8_u1_447_inst:flowthrough inputs: " & " opcode_208 = "& Convert_SLV_To_Hex_String(opcode_208) & " R_BN_446_wire_constant = "& Convert_SLV_To_Hex_String(R_BN_446_wire_constant) & " outputs:" & " EQ_u8_u1_447_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_447_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_447_inst
    process(opcode_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_208, R_BN_446_wire_constant, tmp_var);
      EQ_u8_u1_447_wire <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u32_u32_269_inst flow-through 
    process(LSHR_u32_u32_269_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:LSHR_u32_u32_269_inst:flowthrough inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer) & " outputs:" & " LSHR_u32_u32_269_wire= "  & Convert_SLV_To_Hex_String(LSHR_u32_u32_269_wire));
      --
    end process; 
    -- binary operator LSHR_u32_u32_269_inst
    process(iexec_rd1_final_buffer, iexec_rd2_final_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(iexec_rd1_final_buffer, iexec_rd2_final_buffer, tmp_var);
      LSHR_u32_u32_269_wire <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u32_u32_396_inst flow-through 
    process(bottom_bits_397) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:LSHR_u32_u32_396_inst:flowthrough inputs: " & " is_SRA_385 (guard)= " & Convert_SLV_To_String(is_SRA_385) & " iexec_rd1_final_357_delayed_1_0_388 = "& Convert_SLV_To_Hex_String(iexec_rd1_final_357_delayed_1_0_388) & " iexec_rd2_final_358_delayed_1_0_391 = "& Convert_SLV_To_Hex_String(iexec_rd2_final_358_delayed_1_0_391) & " outputs:" & " bottom_bits_397= "  & Convert_SLV_To_Hex_String(bottom_bits_397));
      --
    end process; 
    -- binary operator LSHR_u32_u32_396_inst
    process(iexec_rd1_final_357_delayed_1_0_388, iexec_rd2_final_358_delayed_1_0_391) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(iexec_rd1_final_357_delayed_1_0_388, iexec_rd2_final_358_delayed_1_0_391, tmp_var);
      bottom_bits_397 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u32_u32_409_inst flow-through 
    process(LSHR_u32_u32_409_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:LSHR_u32_u32_409_inst:flowthrough inputs: " & " is_SRA_385 (guard)= " & Convert_SLV_To_String(is_SRA_385) & " iexec_rd1_final_364_delayed_1_0_400 = "& Convert_SLV_To_Hex_String(iexec_rd1_final_364_delayed_1_0_400) & " R_thirty_one_32_408_wire_constant = "& Convert_SLV_To_Hex_String(R_thirty_one_32_408_wire_constant) & " outputs:" & " LSHR_u32_u32_409_wire= "  & Convert_SLV_To_Hex_String(LSHR_u32_u32_409_wire));
      --
    end process; 
    -- binary operator LSHR_u32_u32_409_inst
    process(iexec_rd1_final_364_delayed_1_0_400) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(iexec_rd1_final_364_delayed_1_0_400, R_thirty_one_32_408_wire_constant, tmp_var);
      LSHR_u32_u32_409_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_434_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NOT_u1_u1_434_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:NOT_u1_u1_434_inst:started:   inputs: " & " is_rs1_neg_431 = "& Convert_SLV_To_Hex_String(is_rs1_neg_431));
          --
        end if; 
        if NOT_u1_u1_434_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:NOT_u1_u1_434_inst:finished:  outputs: " & " NOT_u1_u1_399_399_delayed_1_0_435= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_399_399_delayed_1_0_435));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (32) : NOT_u1_u1_434_inst 
    ApIntNot_group_32: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= is_rs1_neg_431;
      NOT_u1_u1_399_399_delayed_1_0_435 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_434_inst_req_0;
      NOT_u1_u1_434_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_434_inst_req_1;
      NOT_u1_u1_434_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_32_gI: SplitGuardInterface generic map(name => "ApIntNot_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- logger for split-operator OR_u1_u1_450_inst flow-through 
    process(is_Branch_451) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u1_u1_450_inst:flowthrough inputs: " & " AND_u1_u1_444_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_444_wire) & " AND_u1_u1_449_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_449_wire) & " outputs:" & " is_Branch_451= "  & Convert_SLV_To_Hex_String(is_Branch_451));
      --
    end process; 
    -- binary operator OR_u1_u1_450_inst
    process(AND_u1_u1_444_wire, AND_u1_u1_449_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_444_wire, AND_u1_u1_449_wire, tmp_var);
      is_Branch_451 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_233_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if OR_u32_u32_233_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_233_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if OR_u32_u32_233_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_233_inst:finished:  outputs: " & " OR_u32_u32_250_250_delayed_1_0_234= "  & Convert_SLV_To_Hex_String(OR_u32_u32_250_250_delayed_1_0_234));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (34) : OR_u32_u32_233_inst 
    ApIntOr_group_34: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iexec_rd1_final_buffer & iexec_rd2_final_buffer;
      OR_u32_u32_250_250_delayed_1_0_234 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_233_inst_req_0;
      OR_u32_u32_233_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_233_inst_req_1;
      OR_u32_u32_233_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_34_gI: SplitGuardInterface generic map(name => "ApIntOr_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- logger for split-operator OR_u32_u32_285_inst flow-through 
    process(OR_u32_u32_285_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_285_inst:flowthrough inputs: " & " MUX_278_wire = "& Convert_SLV_To_Hex_String(MUX_278_wire) & " MUX_284_wire = "& Convert_SLV_To_Hex_String(MUX_284_wire) & " outputs:" & " OR_u32_u32_285_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_285_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_285_inst
    process(MUX_278_wire, MUX_284_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_278_wire, MUX_284_wire, tmp_var);
      OR_u32_u32_285_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_292_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if OR_u32_u32_292_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_292_inst:started:   inputs: " & " OR_u32_u32_285_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_285_wire) & " MUX_291_wire = "& Convert_SLV_To_Hex_String(MUX_291_wire));
          --
        end if; 
        if OR_u32_u32_292_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_292_inst:finished:  outputs: " & " OR_u32_u32_331_331_delayed_1_0_293= "  & Convert_SLV_To_Hex_String(OR_u32_u32_331_331_delayed_1_0_293));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (36) : OR_u32_u32_292_inst 
    ApIntOr_group_36: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= OR_u32_u32_285_wire & MUX_291_wire;
      OR_u32_u32_331_331_delayed_1_0_293 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_292_inst_req_0;
      OR_u32_u32_292_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_292_inst_req_1;
      OR_u32_u32_292_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_36_gI: SplitGuardInterface generic map(name => "ApIntOr_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- logger for split-operator OR_u32_u32_301_inst flow-through 
    process(OR_u32_u32_301_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_301_inst:flowthrough inputs: " & " AND_u32_u32_230_230_delayed_1_0_239 = "& Convert_SLV_To_Hex_String(AND_u32_u32_230_230_delayed_1_0_239) & " type_cast_300_wire = "& Convert_SLV_To_Hex_String(type_cast_300_wire) & " outputs:" & " OR_u32_u32_301_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_301_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_301_inst
    process(AND_u32_u32_230_230_delayed_1_0_239, type_cast_300_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u32_u32_230_230_delayed_1_0_239, type_cast_300_wire, tmp_var);
      OR_u32_u32_301_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_310_inst flow-through 
    process(OR_u32_u32_310_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_310_inst:flowthrough inputs: " & " MUX_303_wire = "& Convert_SLV_To_Hex_String(MUX_303_wire) & " MUX_309_wire = "& Convert_SLV_To_Hex_String(MUX_309_wire) & " outputs:" & " OR_u32_u32_310_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_310_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_310_inst
    process(MUX_303_wire, MUX_309_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_303_wire, MUX_309_wire, tmp_var);
      OR_u32_u32_310_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_317_inst flow-through 
    process(OR_u32_u32_317_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_317_inst:flowthrough inputs: " & " OR_u32_u32_310_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_310_wire) & " MUX_316_wire = "& Convert_SLV_To_Hex_String(MUX_316_wire) & " outputs:" & " OR_u32_u32_317_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_317_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_317_inst
    process(OR_u32_u32_310_wire, MUX_316_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_310_wire, MUX_316_wire, tmp_var);
      OR_u32_u32_317_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_330_inst flow-through 
    process(OR_u32_u32_330_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_330_inst:flowthrough inputs: " & " MUX_323_wire = "& Convert_SLV_To_Hex_String(MUX_323_wire) & " MUX_329_wire = "& Convert_SLV_To_Hex_String(MUX_329_wire) & " outputs:" & " OR_u32_u32_330_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_330_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_330_inst
    process(MUX_323_wire, MUX_329_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_323_wire, MUX_329_wire, tmp_var);
      OR_u32_u32_330_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_337_inst flow-through 
    process(OR_u32_u32_337_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_337_inst:flowthrough inputs: " & " OR_u32_u32_330_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_330_wire) & " MUX_336_wire = "& Convert_SLV_To_Hex_String(MUX_336_wire) & " outputs:" & " OR_u32_u32_337_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_337_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_337_inst
    process(OR_u32_u32_330_wire, MUX_336_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_330_wire, MUX_336_wire, tmp_var);
      OR_u32_u32_337_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_338_inst flow-through 
    process(OR_u32_u32_338_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_338_inst:flowthrough inputs: " & " OR_u32_u32_317_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_317_wire) & " OR_u32_u32_337_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_337_wire) & " outputs:" & " OR_u32_u32_338_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_338_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_338_inst
    process(OR_u32_u32_317_wire, OR_u32_u32_337_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_317_wire, OR_u32_u32_337_wire, tmp_var);
      OR_u32_u32_338_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_351_inst flow-through 
    process(OR_u32_u32_351_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_351_inst:flowthrough inputs: " & " MUX_344_wire = "& Convert_SLV_To_Hex_String(MUX_344_wire) & " MUX_350_wire = "& Convert_SLV_To_Hex_String(MUX_350_wire) & " outputs:" & " OR_u32_u32_351_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_351_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_351_inst
    process(MUX_344_wire, MUX_350_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_344_wire, MUX_350_wire, tmp_var);
      OR_u32_u32_351_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_358_inst flow-through 
    process(OR_u32_u32_358_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_358_inst:flowthrough inputs: " & " OR_u32_u32_351_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_351_wire) & " MUX_357_wire = "& Convert_SLV_To_Hex_String(MUX_357_wire) & " outputs:" & " OR_u32_u32_358_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_358_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_358_inst
    process(OR_u32_u32_351_wire, MUX_357_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_351_wire, MUX_357_wire, tmp_var);
      OR_u32_u32_358_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_374_inst flow-through 
    process(OR_u32_u32_374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_374_inst:flowthrough inputs: " & " MUX_364_wire = "& Convert_SLV_To_Hex_String(MUX_364_wire) & " MUX_373_wire = "& Convert_SLV_To_Hex_String(MUX_373_wire) & " outputs:" & " OR_u32_u32_374_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_374_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_374_inst
    process(MUX_364_wire, MUX_373_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_364_wire, MUX_373_wire, tmp_var);
      OR_u32_u32_374_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_375_inst flow-through 
    process(OR_u32_u32_375_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_375_inst:flowthrough inputs: " & " OR_u32_u32_358_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_358_wire) & " OR_u32_u32_374_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_374_wire) & " outputs:" & " OR_u32_u32_375_wire= "  & Convert_SLV_To_Hex_String(OR_u32_u32_375_wire));
      --
    end process; 
    -- binary operator OR_u32_u32_375_inst
    process(OR_u32_u32_358_wire, OR_u32_u32_374_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_358_wire, OR_u32_u32_374_wire, tmp_var);
      OR_u32_u32_375_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_376_inst flow-through 
    process(exec_result_initial_377) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_376_inst:flowthrough inputs: " & " OR_u32_u32_338_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_338_wire) & " OR_u32_u32_375_wire = "& Convert_SLV_To_Hex_String(OR_u32_u32_375_wire) & " outputs:" & " exec_result_initial_377= "  & Convert_SLV_To_Hex_String(exec_result_initial_377));
      --
    end process; 
    -- binary operator OR_u32_u32_376_inst
    process(OR_u32_u32_338_wire, OR_u32_u32_375_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_338_wire, OR_u32_u32_375_wire, tmp_var);
      exec_result_initial_377 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u32_u32_420_inst flow-through 
    process(result_for_SRA_421) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:OR_u32_u32_420_inst:flowthrough inputs: " & " is_SRA_385 (guard)= " & Convert_SLV_To_String(is_SRA_385) & " top_bits_415 = "& Convert_SLV_To_Hex_String(top_bits_415) & " bottom_bits_397 = "& Convert_SLV_To_Hex_String(bottom_bits_397) & " outputs:" & " result_for_SRA_421= "  & Convert_SLV_To_Hex_String(result_for_SRA_421));
      --
    end process; 
    -- binary operator OR_u32_u32_420_inst
    process(top_bits_415, bottom_bits_397) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(top_bits_415, bottom_bits_397, tmp_var);
      result_for_SRA_421 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u32_u32_263_inst flow-through 
    process(SHL_u32_u32_263_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:SHL_u32_u32_263_inst:flowthrough inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer) & " outputs:" & " SHL_u32_u32_263_wire= "  & Convert_SLV_To_Hex_String(SHL_u32_u32_263_wire));
      --
    end process; 
    -- binary operator SHL_u32_u32_263_inst
    process(iexec_rd1_final_buffer, iexec_rd2_final_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(iexec_rd1_final_buffer, iexec_rd2_final_buffer, tmp_var);
      SHL_u32_u32_263_wire <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u32_u32_414_inst flow-through 
    process(top_bits_415) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:SHL_u32_u32_414_inst:flowthrough inputs: " & " is_SRA_385 (guard)= " & Convert_SLV_To_String(is_SRA_385) & " SUB_u32_u32_410_wire = "& Convert_SLV_To_Hex_String(SUB_u32_u32_410_wire) & " SUB_u32_u32_413_wire = "& Convert_SLV_To_Hex_String(SUB_u32_u32_413_wire) & " outputs:" & " top_bits_415= "  & Convert_SLV_To_Hex_String(top_bits_415));
      --
    end process; 
    -- binary operator SHL_u32_u32_414_inst
    process(SUB_u32_u32_410_wire, SUB_u32_u32_413_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u32_u32_410_wire, SUB_u32_u32_413_wire, tmp_var);
      top_bits_415 <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u32_u32_258_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if SUB_u32_u32_258_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:SUB_u32_u32_258_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if SUB_u32_u32_258_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:SUB_u32_u32_258_inst:finished:  outputs: " & " SUB_u32_u32_286_286_delayed_1_0_259= "  & Convert_SLV_To_Hex_String(SUB_u32_u32_286_286_delayed_1_0_259));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (51) : SUB_u32_u32_258_inst 
    ApIntSub_group_51: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iexec_rd1_final_buffer & iexec_rd2_final_buffer;
      SUB_u32_u32_286_286_delayed_1_0_259 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_258_inst_req_0;
      SUB_u32_u32_258_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_258_inst_req_1;
      SUB_u32_u32_258_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_51_gI: SplitGuardInterface generic map(name => "ApIntSub_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- logger for split-operator SUB_u32_u32_410_inst flow-through 
    process(SUB_u32_u32_410_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:SUB_u32_u32_410_inst:flowthrough inputs: " & " is_SRA_385 (guard)= " & Convert_SLV_To_String(is_SRA_385) & " R_zero_32_406_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_32_406_wire_constant) & " LSHR_u32_u32_409_wire = "& Convert_SLV_To_Hex_String(LSHR_u32_u32_409_wire) & " outputs:" & " SUB_u32_u32_410_wire= "  & Convert_SLV_To_Hex_String(SUB_u32_u32_410_wire));
      --
    end process; 
    -- binary operator SUB_u32_u32_410_inst
    process(R_zero_32_406_wire_constant, LSHR_u32_u32_409_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_zero_32_406_wire_constant, LSHR_u32_u32_409_wire, tmp_var);
      SUB_u32_u32_410_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u32_u32_413_inst flow-through 
    process(SUB_u32_u32_413_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:SUB_u32_u32_413_inst:flowthrough inputs: " & " is_SRA_385 (guard)= " & Convert_SLV_To_String(is_SRA_385) & " R_thirty_two_32_411_wire_constant = "& Convert_SLV_To_Hex_String(R_thirty_two_32_411_wire_constant) & " iexec_rd2_final_369_delayed_1_0_403 = "& Convert_SLV_To_Hex_String(iexec_rd2_final_369_delayed_1_0_403) & " outputs:" & " SUB_u32_u32_413_wire= "  & Convert_SLV_To_Hex_String(SUB_u32_u32_413_wire));
      --
    end process; 
    -- binary operator SUB_u32_u32_413_inst
    process(R_thirty_two_32_411_wire_constant, iexec_rd2_final_369_delayed_1_0_403) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_thirty_two_32_411_wire_constant, iexec_rd2_final_369_delayed_1_0_403, tmp_var);
      SUB_u32_u32_413_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u32_u1_288_inst flow-through 
    process(UGT_u32_u1_288_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:UGT_u32_u1_288_inst:flowthrough inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer) & " outputs:" & " UGT_u32_u1_288_wire= "  & Convert_SLV_To_Hex_String(UGT_u32_u1_288_wire));
      --
    end process; 
    -- binary operator UGT_u32_u1_288_inst
    process(iexec_rd1_final_buffer, iexec_rd2_final_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(iexec_rd1_final_buffer, iexec_rd2_final_buffer, tmp_var);
      UGT_u32_u1_288_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u32_u1_281_inst flow-through 
    process(ULT_u32_u1_281_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:ULT_u32_u1_281_inst:flowthrough inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer) & " outputs:" & " ULT_u32_u1_281_wire= "  & Convert_SLV_To_Hex_String(ULT_u32_u1_281_wire));
      --
    end process; 
    -- binary operator ULT_u32_u1_281_inst
    process(iexec_rd1_final_buffer, iexec_rd2_final_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(iexec_rd1_final_buffer, iexec_rd2_final_buffer, tmp_var);
      ULT_u32_u1_281_wire <= tmp_var; --
    end process;
    -- logger for split-operator XOR_u32_u32_243_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if XOR_u32_u32_243_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:XOR_u32_u32_243_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if XOR_u32_u32_243_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:XOR_u32_u32_243_inst:finished:  outputs: " & " XOR_u32_u32_259_259_delayed_1_0_244= "  & Convert_SLV_To_Hex_String(XOR_u32_u32_259_259_delayed_1_0_244));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (56) : XOR_u32_u32_243_inst 
    ApIntXnor_group_56: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iexec_rd1_final_buffer & iexec_rd2_final_buffer;
      XOR_u32_u32_259_259_delayed_1_0_244 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_243_inst_req_0;
      XOR_u32_u32_243_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_243_inst_req_1;
      XOR_u32_u32_243_inst_ack_1 <= ackR_unguarded(0);
      ApIntXnor_group_56_gI: SplitGuardInterface generic map(name => "ApIntXnor_group_56_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXnor",
          name => "ApIntXnor_group_56",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- logger for split-operator XOR_u32_u32_248_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if XOR_u32_u32_248_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:XOR_u32_u32_248_inst:started:   inputs: " & " iexec_rd1_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd1_final_buffer) & " iexec_rd2_final_buffer = "& Convert_SLV_To_Hex_String(iexec_rd2_final_buffer));
          --
        end if; 
        if XOR_u32_u32_248_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:iExecStage:DP:XOR_u32_u32_248_inst:finished:  outputs: " & " XOR_u32_u32_267_267_delayed_1_0_249= "  & Convert_SLV_To_Hex_String(XOR_u32_u32_267_267_delayed_1_0_249));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (57) : XOR_u32_u32_248_inst 
    ApIntXor_group_57: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iexec_rd1_final_buffer & iexec_rd2_final_buffer;
      XOR_u32_u32_267_267_delayed_1_0_249 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_248_inst_req_0;
      XOR_u32_u32_248_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_248_inst_req_1;
      XOR_u32_u32_248_inst_ack_1 <= ackR_unguarded(0);
      ApIntXor_group_57_gI: SplitGuardInterface generic map(name => "ApIntXor_group_57_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_57",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- 
  end Block; -- data_path
  -- 
end iExecStage_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity memAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    accessMem_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    accessMem_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    accessMem_request_pipe_read_data : in   std_logic_vector(63 downto 0);
    accessMem_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    accessMem_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    accessMem_response_pipe_write_data : out  std_logic_vector(31 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(42 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(31 downto 0);
    accessMem_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity memAccessDaemon;
architecture memAccessDaemon_arch of memAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal memAccessDaemon_CP_810_start: Boolean;
  signal memAccessDaemon_CP_810_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(9 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_accessMem_request_483_inst_ack_0 : boolean;
  signal do_while_stmt_480_branch_ack_0 : boolean;
  signal RPIPE_accessMem_request_483_inst_ack_1 : boolean;
  signal RPIPE_accessMem_request_483_inst_req_1 : boolean;
  signal call_stmt_501_call_req_1 : boolean;
  signal WPIPE_accessMem_response_502_inst_req_0 : boolean;
  signal WPIPE_accessMem_response_502_inst_ack_0 : boolean;
  signal do_while_stmt_480_branch_req_0 : boolean;
  signal call_stmt_501_call_ack_1 : boolean;
  signal WPIPE_accessMem_response_502_inst_ack_1 : boolean;
  signal RPIPE_accessMem_request_483_inst_req_0 : boolean;
  signal do_while_stmt_480_branch_ack_1 : boolean;
  signal WPIPE_accessMem_response_502_inst_req_1 : boolean;
  signal call_stmt_501_call_ack_0 : boolean;
  signal call_stmt_501_call_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "memAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  memAccessDaemon_CP_810_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "memAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memAccessDaemon_CP_810_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= memAccessDaemon_CP_810_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memAccessDaemon_CP_810_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,memAccessDaemon_CP_810_start,"memAccessDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,memAccessDaemon_CP_810_symbol, "memAccessDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  memAccessDaemon_CP_810: Block -- control-path 
    signal memAccessDaemon_CP_810_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    memAccessDaemon_CP_810_elements(0) <= memAccessDaemon_CP_810_start;
    memAccessDaemon_CP_810_symbol <= memAccessDaemon_CP_810_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_479/$entry
      -- CP-element group 0: 	 branch_block_stmt_479/do_while_stmt_480__entry__
      -- CP-element group 0: 	 branch_block_stmt_479/branch_block_stmt_479__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	24 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_479/do_while_stmt_480__exit__
      -- CP-element group 1: 	 branch_block_stmt_479/$exit
      -- CP-element group 1: 	 branch_block_stmt_479/branch_block_stmt_479__exit__
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_810_elements(1) <= memAccessDaemon_CP_810_elements(24);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480__entry__
      -- CP-element group 2: 	 branch_block_stmt_479/do_while_stmt_480/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_810_elements(2) <= memAccessDaemon_CP_810_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	24 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480__exit__
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon_CP_810_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_479/do_while_stmt_480/loop_back
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon_CP_810_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	21 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	22 
    -- CP-element group 5: 	23 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_479/do_while_stmt_480/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_479/do_while_stmt_480/condition_done
      -- CP-element group 5: 	 branch_block_stmt_479/do_while_stmt_480/loop_taken/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_810_elements(5) <= memAccessDaemon_CP_810_elements(21);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	20 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_479/do_while_stmt_480/loop_body_done
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_810_elements(6) <= memAccessDaemon_CP_810_elements(20);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_810_elements(7) <= memAccessDaemon_CP_810_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_810_elements(8) <= memAccessDaemon_CP_810_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	21 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon_CP_810_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_sample_start_
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_accessMem_request_483_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_810_elements(10), ack => RPIPE_accessMem_request_483_inst_req_0); -- 
    memAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_810_elements(9) & memAccessDaemon_CP_810_elements(13);
      gj_memAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_810_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_update_start_
      -- CP-element group 11: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Update/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_accessMem_request_483_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_810_elements(11), ack => RPIPE_accessMem_request_483_inst_req_1); -- 
    memAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_810_elements(12) & memAccessDaemon_CP_810_elements(16);
      gj_memAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_810_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_sample_completed_
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_accessMem_request_483_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_accessMem_request_483_inst_ack_0, ack => memAccessDaemon_CP_810_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/RPIPE_accessMem_request_483_Update/$exit
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_accessMem_request_483_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_accessMem_request_483_inst_ack_1, ack => memAccessDaemon_CP_810_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Sample/crr
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_501_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_810_elements(14), ack => call_stmt_501_call_req_0); -- 
    memAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_810_elements(13) & memAccessDaemon_CP_810_elements(16);
      gj_memAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_810_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_update_start_
      -- CP-element group 15: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Update/ccr
      -- CP-element group 15: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Update/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_501_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_810_elements(15), ack => call_stmt_501_call_req_1); -- 
    memAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memAccessDaemon_CP_810_elements(19);
      gj_memAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_810_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Sample/cra
      -- CP-element group 16: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Sample/$exit
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_501_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_501_call_ack_0, ack => memAccessDaemon_CP_810_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Update/cca
      -- CP-element group 17: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/call_stmt_501_Update/$exit
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_501_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_501_call_ack_1, ack => memAccessDaemon_CP_810_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Sample/req
      -- CP-element group 18: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Sample/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_accessMem_response_502_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_810_elements(18), ack => WPIPE_accessMem_response_502_inst_req_0); -- 
    memAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_810_elements(17) & memAccessDaemon_CP_810_elements(20);
      gj_memAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_810_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Sample/ack
      -- CP-element group 19: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Update/req
      -- CP-element group 19: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_update_start_
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_accessMem_response_502_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_accessMem_response_502_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accessMem_response_502_inst_ack_0, ack => memAccessDaemon_CP_810_elements(19)); -- 
    req_876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_810_elements(19), ack => WPIPE_accessMem_response_502_inst_req_1); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (4) 
      -- CP-element group 20: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/$exit
      -- CP-element group 20: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_Update/ack
      -- CP-element group 20: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/WPIPE_accessMem_response_502_update_completed_
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_accessMem_response_502_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accessMem_response_502_inst_ack_1, ack => memAccessDaemon_CP_810_elements(20)); -- 
    -- CP-element group 21:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	5 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/condition_evaluated
      -- CP-element group 21: 	 branch_block_stmt_479/do_while_stmt_480/do_while_stmt_480_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:do_while_stmt_480_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_810_elements(21), ack => do_while_stmt_480_branch_req_0); -- 
    -- Element group memAccessDaemon_CP_810_elements(21) is a control-delay.
    cp_element_21_delay: control_delay_element  generic map(name => " 21_delay", delay_value => 1)  port map(req => memAccessDaemon_CP_810_elements(9), ack => memAccessDaemon_CP_810_elements(21), clk => clk, reset =>reset);
    -- CP-element group 22:  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_479/do_while_stmt_480/loop_exit/$exit
      -- CP-element group 22: 	 branch_block_stmt_479/do_while_stmt_480/loop_exit/ack
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:do_while_stmt_480_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_480_branch_ack_0, ack => memAccessDaemon_CP_810_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	5 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_479/do_while_stmt_480/loop_taken/$exit
      -- CP-element group 23: 	 branch_block_stmt_479/do_while_stmt_480/loop_taken/ack
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:do_while_stmt_480_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_480_branch_ack_1, ack => memAccessDaemon_CP_810_elements(23)); -- 
    -- CP-element group 24:  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	3 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	1 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_479/do_while_stmt_480/$exit
      -- 
    -- logger for CP element group memAccessDaemon_CP_810_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_810_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_810_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_810_elements(24) <= memAccessDaemon_CP_810_elements(3);
    memAccessDaemon_do_while_stmt_480_terminator_887: loop_terminator -- 
      generic map (name => " memAccessDaemon_do_while_stmt_480_terminator_887", max_iterations_in_flight =>20) 
      port map(loop_body_exit => memAccessDaemon_CP_810_elements(6),loop_continue => memAccessDaemon_CP_810_elements(23),loop_terminate => memAccessDaemon_CP_810_elements(22),loop_back => memAccessDaemon_CP_810_elements(4),loop_exit => memAccessDaemon_CP_810_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_835_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= memAccessDaemon_CP_810_elements(7);
        preds(1)  <= memAccessDaemon_CP_810_elements(8);
        entry_tmerge_835 : transition_merge -- 
          generic map(name => " entry_tmerge_835")
          port map (preds => preds, symbol_out => memAccessDaemon_CP_810_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addr_492 : std_logic_vector(9 downto 0);
    signal cmd_1_484 : std_logic_vector(63 downto 0);
    signal konst_506_wire_constant : std_logic_vector(0 downto 0);
    signal rdata_501 : std_logic_vector(31 downto 0);
    signal rwbar_496 : std_logic_vector(0 downto 0);
    signal wdata_488 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_506_wire_constant <= "1";
    -- logger for split-operator slice_487_inst flow-through 
    process(wdata_488) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:slice_487_inst:flowthrough inputs: " & " cmd_1_484 = "& Convert_SLV_To_Hex_String(cmd_1_484) & " outputs:" & " wdata_488= "  & Convert_SLV_To_Hex_String(wdata_488));
      --
    end process; 
    -- flow-through slice operator slice_487_inst
    wdata_488 <= cmd_1_484(63 downto 32);
    -- logger for split-operator slice_491_inst flow-through 
    process(addr_492) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:slice_491_inst:flowthrough inputs: " & " cmd_1_484 = "& Convert_SLV_To_Hex_String(cmd_1_484) & " outputs:" & " addr_492= "  & Convert_SLV_To_Hex_String(addr_492));
      --
    end process; 
    -- flow-through slice operator slice_491_inst
    addr_492 <= cmd_1_484(31 downto 22);
    -- logger for split-operator slice_495_inst flow-through 
    process(rwbar_496) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:slice_495_inst:flowthrough inputs: " & " cmd_1_484 = "& Convert_SLV_To_Hex_String(cmd_1_484) & " outputs:" & " rwbar_496= "  & Convert_SLV_To_Hex_String(rwbar_496));
      --
    end process; 
    -- flow-through slice operator slice_495_inst
    rwbar_496 <= cmd_1_484(0 downto 0);
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_480_branch_req_0," req0 do_while_stmt_480_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_480_branch_ack_0," ack0 do_while_stmt_480_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_480_branch_ack_1," ack1 do_while_stmt_480_branch");
    do_while_stmt_480_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_506_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_480_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_480_branch_req_0,
          ack0 => do_while_stmt_480_branch_ack_0,
          ack1 => do_while_stmt_480_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_accessMem_request_483_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_accessMem_request_483_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:RPIPE_accessMem_request_483_inst:started:   PipeRead from accessMem_request inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_accessMem_request_483_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:RPIPE_accessMem_request_483_inst:finished:  outputs: " & " cmd_1_484= "  & Convert_SLV_To_Hex_String(cmd_1_484));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_accessMem_request_483_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_accessMem_request_483_inst_req_0;
      RPIPE_accessMem_request_483_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_accessMem_request_483_inst_req_1;
      RPIPE_accessMem_request_483_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      cmd_1_484 <= data_out(63 downto 0);
      accessMem_request_read_0_gI: SplitGuardInterface generic map(name => "accessMem_request_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      accessMem_request_read_0: InputPortRevised -- 
        generic map ( name => "accessMem_request_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => accessMem_request_pipe_read_req(0),
          oack => accessMem_request_pipe_read_ack(0),
          odata => accessMem_request_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_accessMem_response_502_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_accessMem_response_502_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:WPIPE_accessMem_response_502_inst:started:   PipeWrite to accessMem_response inputs: " & " rdata_501 = "& Convert_SLV_To_Hex_String(rdata_501));
          --
        end if; 
        if WPIPE_accessMem_response_502_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:WPIPE_accessMem_response_502_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_accessMem_response_502_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_accessMem_response_502_inst_req_0;
      WPIPE_accessMem_response_502_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_accessMem_response_502_inst_req_1;
      WPIPE_accessMem_response_502_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= rdata_501;
      accessMem_response_write_0_gI: SplitGuardInterface generic map(name => "accessMem_response_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      accessMem_response_write_0: OutputPortRevised -- 
        generic map ( name => "accessMem_response", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => accessMem_response_pipe_write_req(0),
          oack => accessMem_response_pipe_write_ack(0),
          odata => accessMem_response_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_501_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_501_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:call_stmt_501_call:started:  Call to module accessMem inputs: " & " rwbar_496 = "& Convert_SLV_To_Hex_String(rwbar_496) & " addr_492 = "& Convert_SLV_To_Hex_String(addr_492) & " wdata_488 = "& Convert_SLV_To_Hex_String(wdata_488));
          --
        end if; 
        if call_stmt_501_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:call_stmt_501_call:finished:  outputs: " & " rdata_501= "  & Convert_SLV_To_Hex_String(rdata_501));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_501_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 7);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_501_call_req_0;
      call_stmt_501_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_501_call_req_1;
      call_stmt_501_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rwbar_496 & addr_492 & wdata_488;
      rdata_501 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(42 downto 0),
          tagR => accessMem_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(31 downto 0),
          tagL => accessMem_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end memAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity processor_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_processor_pipe_read_req : out  std_logic_vector(0 downto 0);
    start_processor_pipe_read_ack : in   std_logic_vector(0 downto 0);
    start_processor_pipe_read_data : in   std_logic_vector(7 downto 0);
    processor_result_pipe_write_req : out  std_logic_vector(0 downto 0);
    processor_result_pipe_write_ack : in   std_logic_vector(0 downto 0);
    processor_result_pipe_write_data : out  std_logic_vector(31 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(42 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(31 downto 0);
    accessMem_return_tag :  in   std_logic_vector(1 downto 0);
    iExecStage_call_reqs : out  std_logic_vector(0 downto 0);
    iExecStage_call_acks : in   std_logic_vector(0 downto 0);
    iExecStage_call_data : out  std_logic_vector(169 downto 0);
    iExecStage_call_tag  :  out  std_logic_vector(0 downto 0);
    iExecStage_return_reqs : out  std_logic_vector(0 downto 0);
    iExecStage_return_acks : in   std_logic_vector(0 downto 0);
    iExecStage_return_data : in   std_logic_vector(138 downto 0);
    iExecStage_return_tag :  in   std_logic_vector(0 downto 0);
    accessReg_call_reqs : out  std_logic_vector(0 downto 0);
    accessReg_call_acks : in   std_logic_vector(0 downto 0);
    accessReg_call_data : out  std_logic_vector(58 downto 0);
    accessReg_call_tag  :  out  std_logic_vector(0 downto 0);
    accessReg_return_reqs : out  std_logic_vector(0 downto 0);
    accessReg_return_acks : in   std_logic_vector(0 downto 0);
    accessReg_return_data : in   std_logic_vector(63 downto 0);
    accessReg_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity processor_daemon;
architecture processor_daemon_arch of processor_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal processor_daemon_CP_891_start: Boolean;
  signal processor_daemon_CP_891_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(9 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component iExecStage is -- 
    generic (tag_length : integer); 
    port ( -- 
      iexec_state : in  std_logic_vector(105 downto 0);
      iexec_rd1_final : in  std_logic_vector(31 downto 0);
      iexec_rd2_final : in  std_logic_vector(31 downto 0);
      next_dcache_state : out  std_logic_vector(138 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessReg is -- 
    generic (tag_length : integer); 
    port ( -- 
      valid_1 : in  std_logic_vector(0 downto 0);
      addr_1 : in  std_logic_vector(7 downto 0);
      valid_2 : in  std_logic_vector(0 downto 0);
      addr_2 : in  std_logic_vector(7 downto 0);
      valid_w : in  std_logic_vector(0 downto 0);
      addr_w : in  std_logic_vector(7 downto 0);
      data_to_be_written : in  std_logic_vector(31 downto 0);
      read_data_1 : out  std_logic_vector(31 downto 0);
      read_data_2 : out  std_logic_vector(31 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component scoreBoard_Volatile is -- 
    port ( -- 
      clk, reset: in std_logic; 
      ifetch_state : in  std_logic_vector(9 downto 0);
      icache_state : in  std_logic_vector(9 downto 0);
      idecode_state : in  std_logic_vector(41 downto 0);
      iregfile_state : in  std_logic_vector(41 downto 0);
      iexec_state : in  std_logic_vector(105 downto 0);
      dcache_state : in  std_logic_vector(138 downto 0);
      iretire_state : in  std_logic_vector(138 downto 0);
      ifetch_actions : out  std_logic_vector(9 downto 0);
      icache_actions : out  std_logic_vector(9 downto 0);
      idecode_actions : out  std_logic_vector(41 downto 0);
      iregfile_actions : out  std_logic_vector(4 downto 0);
      iexec_actions : out  std_logic_vector(3 downto 0);
      dcache_actions : out  std_logic_vector(2 downto 0);
      ex_Unconditional_JUMP : out  std_logic_vector(0 downto 0);
      is_Branch_Hazard : out  std_logic_vector(0 downto 0);
      flush_ifetch : out  std_logic_vector(0 downto 0);
      flush_icache : out  std_logic_vector(0 downto 0);
      flush_idecode : out  std_logic_vector(0 downto 0);
      flush_reg : out  std_logic_vector(0 downto 0);
      flush_iexec : out  std_logic_vector(0 downto 0);
      flush_dcache : out  std_logic_vector(0 downto 0);
      stall_first_4 : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal phi_stmt_933_req_1 : boolean;
  signal if_stmt_926_branch_ack_0 : boolean;
  signal RPIPE_start_processor_924_inst_req_0 : boolean;
  signal RPIPE_start_processor_924_inst_req_1 : boolean;
  signal RPIPE_start_processor_924_inst_ack_0 : boolean;
  signal W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_0 : boolean;
  signal if_stmt_926_branch_req_0 : boolean;
  signal MUX_1141_inst_ack_0 : boolean;
  signal next_ifetch_state_1358_936_buf_ack_0 : boolean;
  signal W_flush_dcache_1221_delayed_4_0_1134_inst_req_0 : boolean;
  signal phi_stmt_937_req_1 : boolean;
  signal next_ifetch_state_1358_936_buf_req_0 : boolean;
  signal phi_stmt_933_req_0 : boolean;
  signal phi_stmt_933_ack_0 : boolean;
  signal W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_0 : boolean;
  signal call_stmt_1133_call_ack_0 : boolean;
  signal phi_stmt_945_req_1 : boolean;
  signal W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_0 : boolean;
  signal MUX_1141_inst_ack_1 : boolean;
  signal call_stmt_1133_call_req_0 : boolean;
  signal do_while_stmt_931_branch_req_0 : boolean;
  signal phi_stmt_937_ack_0 : boolean;
  signal next_ifetch_state_1358_936_buf_req_1 : boolean;
  signal RPIPE_start_processor_924_inst_ack_1 : boolean;
  signal phi_stmt_937_req_0 : boolean;
  signal next_ifetch_state_1358_936_buf_ack_1 : boolean;
  signal W_flush_dcache_1221_delayed_4_0_1134_inst_ack_0 : boolean;
  signal if_stmt_926_branch_ack_1 : boolean;
  signal call_stmt_1175_call_ack_0 : boolean;
  signal CONCAT_u24_u64_1299_inst_ack_1 : boolean;
  signal n_icache_state_998_940_buf_ack_1 : boolean;
  signal n_icache_state_998_940_buf_req_1 : boolean;
  signal MUX_1141_inst_req_1 : boolean;
  signal n_icache_state_998_940_buf_ack_0 : boolean;
  signal n_idecode_state_1021_944_buf_ack_1 : boolean;
  signal n_idecode_state_1021_944_buf_req_1 : boolean;
  signal n_idecode_state_1021_944_buf_ack_0 : boolean;
  signal n_idecode_state_1021_944_buf_req_0 : boolean;
  signal n_icache_state_998_940_buf_req_0 : boolean;
  signal CONCAT_u16_u32_1259_inst_ack_0 : boolean;
  signal W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_1 : boolean;
  signal phi_stmt_941_ack_0 : boolean;
  signal phi_stmt_941_req_0 : boolean;
  signal W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_1 : boolean;
  signal phi_stmt_941_req_1 : boolean;
  signal W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_1 : boolean;
  signal MUX_1141_inst_req_0 : boolean;
  signal WPIPE_processor_result_1370_inst_ack_1 : boolean;
  signal W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_1 : boolean;
  signal CONCAT_u16_u32_1259_inst_ack_1 : boolean;
  signal WPIPE_processor_result_1370_inst_ack_0 : boolean;
  signal W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_1 : boolean;
  signal call_stmt_1133_call_req_1 : boolean;
  signal W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_1 : boolean;
  signal W_iregfile_pc_1342_delayed_7_0_1261_inst_req_0 : boolean;
  signal call_stmt_1133_call_ack_1 : boolean;
  signal W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_1 : boolean;
  signal call_stmt_1175_call_req_1 : boolean;
  signal call_stmt_1175_call_ack_1 : boolean;
  signal W_flush_dcache_1221_delayed_4_0_1134_inst_req_1 : boolean;
  signal CONCAT_u16_u32_1259_inst_req_1 : boolean;
  signal W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_0 : boolean;
  signal W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_0 : boolean;
  signal call_stmt_1175_call_req_0 : boolean;
  signal W_flush_dcache_1221_delayed_4_0_1134_inst_ack_1 : boolean;
  signal phi_stmt_945_req_0 : boolean;
  signal W_flush_iexec_1330_delayed_7_0_1249_inst_ack_1 : boolean;
  signal do_while_stmt_931_branch_ack_1 : boolean;
  signal phi_stmt_945_ack_0 : boolean;
  signal WPIPE_processor_result_1370_inst_req_1 : boolean;
  signal W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_1 : boolean;
  signal CONCAT_u24_u64_1299_inst_ack_0 : boolean;
  signal CONCAT_u24_u64_1299_inst_req_0 : boolean;
  signal n_iregfile_state_1030_948_buf_req_0 : boolean;
  signal n_iregfile_state_1030_948_buf_ack_0 : boolean;
  signal W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_0 : boolean;
  signal n_iregfile_state_1030_948_buf_req_1 : boolean;
  signal n_iregfile_state_1030_948_buf_ack_1 : boolean;
  signal CONCAT_u1_u11_1307_inst_ack_0 : boolean;
  signal W_flush_iexec_1330_delayed_7_0_1249_inst_req_1 : boolean;
  signal W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_0 : boolean;
  signal phi_stmt_949_req_1 : boolean;
  signal W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_0 : boolean;
  signal phi_stmt_949_req_0 : boolean;
  signal phi_stmt_949_ack_0 : boolean;
  signal W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_1 : boolean;
  signal W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_1 : boolean;
  signal W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_0 : boolean;
  signal n_iexec_state_1275_952_buf_req_0 : boolean;
  signal n_iexec_state_1275_952_buf_ack_0 : boolean;
  signal CONCAT_u1_u11_1307_inst_req_0 : boolean;
  signal n_iexec_state_1275_952_buf_req_1 : boolean;
  signal n_iexec_state_1275_952_buf_ack_1 : boolean;
  signal phi_stmt_953_req_1 : boolean;
  signal W_flush_iexec_1330_delayed_7_0_1249_inst_ack_0 : boolean;
  signal phi_stmt_953_req_0 : boolean;
  signal W_flush_iexec_1330_delayed_7_0_1249_inst_req_0 : boolean;
  signal do_while_stmt_931_branch_ack_0 : boolean;
  signal phi_stmt_953_ack_0 : boolean;
  signal W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_0 : boolean;
  signal CONCAT_u1_u11_1307_inst_ack_1 : boolean;
  signal W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_0 : boolean;
  signal n_dcache_state_1142_956_buf_req_0 : boolean;
  signal n_dcache_state_1142_956_buf_ack_0 : boolean;
  signal n_dcache_state_1142_956_buf_req_1 : boolean;
  signal n_dcache_state_1142_956_buf_ack_1 : boolean;
  signal phi_stmt_957_req_1 : boolean;
  signal phi_stmt_957_req_0 : boolean;
  signal phi_stmt_957_ack_0 : boolean;
  signal CONCAT_u1_u11_1307_inst_req_1 : boolean;
  signal EQ_u8_u1_1279_inst_ack_1 : boolean;
  signal EQ_u8_u1_1279_inst_req_1 : boolean;
  signal n_iRetire_state_1317_960_buf_req_0 : boolean;
  signal n_iRetire_state_1317_960_buf_ack_0 : boolean;
  signal W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_1 : boolean;
  signal W_dcache_rd2_1365_delayed_7_0_1301_inst_req_1 : boolean;
  signal n_iRetire_state_1317_960_buf_req_1 : boolean;
  signal n_iRetire_state_1317_960_buf_ack_1 : boolean;
  signal call_stmt_989_call_req_0 : boolean;
  signal call_stmt_989_call_ack_0 : boolean;
  signal call_stmt_1224_call_ack_1 : boolean;
  signal call_stmt_989_call_req_1 : boolean;
  signal call_stmt_989_call_ack_1 : boolean;
  signal EQ_u8_u1_1279_inst_ack_0 : boolean;
  signal EQ_u8_u1_1279_inst_req_0 : boolean;
  signal call_stmt_1224_call_req_1 : boolean;
  signal W_flush_idecode_1058_delayed_7_0_999_inst_req_0 : boolean;
  signal W_flush_idecode_1058_delayed_7_0_999_inst_ack_0 : boolean;
  signal W_flush_idecode_1058_delayed_7_0_999_inst_req_1 : boolean;
  signal W_flush_idecode_1058_delayed_7_0_999_inst_ack_1 : boolean;
  signal W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_0 : boolean;
  signal CONCAT_u24_u64_1299_inst_req_1 : boolean;
  signal WPIPE_processor_result_1370_inst_req_0 : boolean;
  signal W_dcache_rd2_1365_delayed_7_0_1301_inst_req_0 : boolean;
  signal W_stall_first_4_1060_delayed_7_0_1002_inst_req_0 : boolean;
  signal W_stall_first_4_1060_delayed_7_0_1002_inst_ack_0 : boolean;
  signal call_stmt_1224_call_ack_0 : boolean;
  signal W_stall_first_4_1060_delayed_7_0_1002_inst_req_1 : boolean;
  signal W_stall_first_4_1060_delayed_7_0_1002_inst_ack_1 : boolean;
  signal W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_1 : boolean;
  signal CONCAT_u16_u32_1259_inst_req_0 : boolean;
  signal call_stmt_1224_call_req_0 : boolean;
  signal W_idecode_state_1061_delayed_7_0_1005_inst_req_0 : boolean;
  signal W_idecode_state_1061_delayed_7_0_1005_inst_ack_0 : boolean;
  signal W_idecode_state_1061_delayed_7_0_1005_inst_req_1 : boolean;
  signal W_idecode_state_1061_delayed_7_0_1005_inst_ack_1 : boolean;
  signal W_iregfile_pc_1342_delayed_7_0_1261_inst_req_1 : boolean;
  signal W_icache_state_1063_delayed_7_0_1008_inst_req_0 : boolean;
  signal W_icache_state_1063_delayed_7_0_1008_inst_ack_0 : boolean;
  signal W_icache_state_1063_delayed_7_0_1008_inst_req_1 : boolean;
  signal W_icache_state_1063_delayed_7_0_1008_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "processor_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  processor_daemon_CP_891_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "processor_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= processor_daemon_CP_891_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= processor_daemon_CP_891_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= processor_daemon_CP_891_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,processor_daemon_CP_891_start,"processor_daemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,processor_daemon_CP_891_symbol, "processor_daemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  processor_daemon_CP_891: Block -- control-path 
    signal processor_daemon_CP_891_elements: BooleanArray(247 downto 0);
    -- 
  begin -- 
    processor_daemon_CP_891_elements(0) <= processor_daemon_CP_891_start;
    processor_daemon_CP_891_symbol <= processor_daemon_CP_891_elements(4);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	247 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_921/$entry
      -- CP-element group 0: 	 branch_block_stmt_921/branch_block_stmt_921__entry__
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922__entry__
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922__entry___PhiReq/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	247 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:RPIPE_start_processor_924_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:RPIPE_start_processor_924_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_start_processor_924_inst_ack_0, ack => processor_daemon_CP_891_elements(1)); -- 
    cr_920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(1), ack => RPIPE_start_processor_924_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926__entry__
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_else_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Update/ca
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/branch_req
      -- CP-element group 2: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/EQ_u8_u1_929_place
      -- CP-element group 2: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/EQ_u8_u1_929_inputs/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/SplitProtocol/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/assign_stmt_925__exit__
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_eval_test/EQ_u8_u1_929/EQ_u8_u1_929_inputs/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_926_if_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/assign_stmt_925/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:RPIPE_start_processor_924_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:if_stmt_926_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_start_processor_924_inst_ack_1, ack => processor_daemon_CP_891_elements(2)); -- 
    branch_req_948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(2), ack => if_stmt_926_branch_req_0); -- 
    -- CP-element group 3:  transition  place  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_921/branch_block_stmt_930/branch_block_stmt_930__entry__
      -- CP-element group 3: 	 branch_block_stmt_921/branch_block_stmt_930/$entry
      -- CP-element group 3: 	 branch_block_stmt_921/if_stmt_926_if_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_921/branch_block_stmt_930__entry__
      -- CP-element group 3: 	 branch_block_stmt_921/if_stmt_926_if_link/if_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931__entry__
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:if_stmt_926_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_926_branch_ack_1, ack => processor_daemon_CP_891_elements(3)); -- 
    -- CP-element group 4:  merge  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_921/if_stmt_926_else_link/else_choice_transition
      -- CP-element group 4: 	 branch_block_stmt_921/if_stmt_926_else_link/$exit
      -- CP-element group 4: 	 branch_block_stmt_921/if_stmt_926__exit__
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 branch_block_stmt_921/branch_block_stmt_921__exit__
      -- CP-element group 4: 	 branch_block_stmt_921/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:if_stmt_926_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_926_branch_ack_0, ack => processor_daemon_CP_891_elements(4)); -- 
    -- CP-element group 5:  transition  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	246 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	247 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 branch_block_stmt_921/branch_block_stmt_930/$exit
      -- CP-element group 5: 	 branch_block_stmt_921/check_for_start
      -- CP-element group 5: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931__exit__
      -- CP-element group 5: 	 branch_block_stmt_921/branch_block_stmt_930/branch_block_stmt_930__exit__
      -- CP-element group 5: 	 branch_block_stmt_921/branch_block_stmt_930__exit__
      -- CP-element group 5: 	 branch_block_stmt_921/check_for_start_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_921/check_for_start_PhiReq/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(5) <= processor_daemon_CP_891_elements(246);
    -- CP-element group 6:  transition  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	12 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931__entry__
      -- CP-element group 6: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(6) <= processor_daemon_CP_891_elements(3);
    -- CP-element group 7:  merge  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	246 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931__exit__
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(7) is bound as output of CP function.
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_back
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(8) is bound as output of CP function.
    -- CP-element group 9:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	244 
    -- CP-element group 9: 	245 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/condition_done
      -- CP-element group 9: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_taken/$entry
      -- CP-element group 9: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_exit/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(9) <= processor_daemon_CP_891_elements(14);
    -- CP-element group 10:  branch  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	243 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_body_done
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(10) <= processor_daemon_CP_891_elements(243);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	120 
    -- CP-element group 11: 	25 
    -- CP-element group 11: 	44 
    -- CP-element group 11: 	63 
    -- CP-element group 11: 	82 
    -- CP-element group 11: 	101 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(11) <= processor_daemon_CP_891_elements(8);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	6 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	122 
    -- CP-element group 12: 	27 
    -- CP-element group 12: 	46 
    -- CP-element group 12: 	65 
    -- CP-element group 12: 	84 
    -- CP-element group 12: 	103 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(12) <= processor_daemon_CP_891_elements(6);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	133 
    -- CP-element group 13: 	134 
    -- CP-element group 13: 	241 
    -- CP-element group 13: 	114 
    -- CP-element group 13: 	115 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	20 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	39 
    -- CP-element group 13: 	57 
    -- CP-element group 13: 	58 
    -- CP-element group 13: 	76 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	95 
    -- CP-element group 13: 	96 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/$entry
      -- CP-element group 13: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/loop_body_start
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(13) is bound as output of CP function.
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	241 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/condition_evaluated
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:do_while_stmt_931_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(14), ack => do_while_stmt_931_branch_req_0); -- 
    processor_daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(241) & processor_daemon_CP_891_elements(18);
      gj_processor_daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	133 
    -- CP-element group 15: 	114 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	57 
    -- CP-element group 15: 	76 
    -- CP-element group 15: 	95 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	116 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	40 
    -- CP-element group 15: 	59 
    -- CP-element group 15: 	78 
    -- CP-element group 15: 	97 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/aggregated_phi_sample_req
      -- CP-element group 15: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(133) & processor_daemon_CP_891_elements(114) & processor_daemon_CP_891_elements(19) & processor_daemon_CP_891_elements(38) & processor_daemon_CP_891_elements(57) & processor_daemon_CP_891_elements(76) & processor_daemon_CP_891_elements(95) & processor_daemon_CP_891_elements(18);
      gj_processor_daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	135 
    -- CP-element group 16: 	117 
    -- CP-element group 16: 	22 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	79 
    -- CP-element group 16: 	98 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	243 
    -- CP-element group 16: 	195 
    -- CP-element group 16: 	199 
    -- CP-element group 16: 	203 
    -- CP-element group 16: 	179 
    -- CP-element group 16: 	227 
    -- CP-element group 16: 	231 
    -- CP-element group 16: 	235 
    -- CP-element group 16: 	207 
    -- CP-element group 16: 	211 
    -- CP-element group 16: 	215 
    -- CP-element group 16: 	219 
    -- CP-element group 16: 	223 
    -- CP-element group 16: 	159 
    -- CP-element group 16: 	163 
    -- CP-element group 16: 	167 
    -- CP-element group 16: 	151 
    -- CP-element group 16: 	155 
    -- CP-element group 16: 	183 
    -- CP-element group 16: 	187 
    -- CP-element group 16: 	191 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	133 
    -- CP-element group 16: 	114 
    -- CP-element group 16: 	19 
    -- CP-element group 16: 	38 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	76 
    -- CP-element group 16: 	95 
    -- CP-element group 16:  members (8) 
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/aggregated_phi_sample_ack
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(135) & processor_daemon_CP_891_elements(117) & processor_daemon_CP_891_elements(22) & processor_daemon_CP_891_elements(41) & processor_daemon_CP_891_elements(60) & processor_daemon_CP_891_elements(79) & processor_daemon_CP_891_elements(98);
      gj_processor_daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	134 
    -- CP-element group 17: 	115 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	39 
    -- CP-element group 17: 	58 
    -- CP-element group 17: 	77 
    -- CP-element group 17: 	96 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	118 
    -- CP-element group 17: 	23 
    -- CP-element group 17: 	42 
    -- CP-element group 17: 	61 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	99 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/aggregated_phi_update_req
      -- CP-element group 17: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(134) & processor_daemon_CP_891_elements(115) & processor_daemon_CP_891_elements(20) & processor_daemon_CP_891_elements(39) & processor_daemon_CP_891_elements(58) & processor_daemon_CP_891_elements(77) & processor_daemon_CP_891_elements(96);
      gj_processor_daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	136 
    -- CP-element group 18: 	119 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	81 
    -- CP-element group 18: 	100 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100);
      gj_processor_daemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	16 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(16);
      gj_processor_daemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	13 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	200 
    -- CP-element group 20: 	172 
    -- CP-element group 20: 	176 
    -- CP-element group 20: 	208 
    -- CP-element group 20: 	160 
    -- CP-element group 20: 	156 
    -- CP-element group 20: 	184 
    -- CP-element group 20: 	188 
    -- CP-element group 20: 	192 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(200) & processor_daemon_CP_891_elements(172) & processor_daemon_CP_891_elements(176) & processor_daemon_CP_891_elements(208) & processor_daemon_CP_891_elements(160) & processor_daemon_CP_891_elements(156) & processor_daemon_CP_891_elements(184) & processor_daemon_CP_891_elements(188) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(21) <= processor_daemon_CP_891_elements(15);
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	16 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(23) <= processor_daemon_CP_891_elements(17);
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	198 
    -- CP-element group 24: 	170 
    -- CP-element group 24: 	174 
    -- CP-element group 24: 	206 
    -- CP-element group 24: 	154 
    -- CP-element group 24: 	158 
    -- CP-element group 24: 	182 
    -- CP-element group 24: 	186 
    -- CP-element group 24: 	190 
    -- CP-element group 24: 	18 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	11 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_loopback_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(25) <= processor_daemon_CP_891_elements(11);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_loopback_sample_req
      -- CP-element group 26: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_loopback_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_933_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_933_loopback_sample_req_997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_933_loopback_sample_req_997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(26), ack => phi_stmt_933_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	12 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_entry_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(27) <= processor_daemon_CP_891_elements(12);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_entry_sample_req
      -- CP-element group 28: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_entry_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_933_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_933_entry_sample_req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_933_entry_sample_req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(28), ack => phi_stmt_933_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_phi_mux_ack
      -- CP-element group 29: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_933_phi_mux_ack_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_933_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_933_phi_mux_ack_1003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_933_ack_0, ack => processor_daemon_CP_891_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(32) <= processor_daemon_CP_891_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_one_10_935_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(33) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(31), ack => processor_daemon_CP_891_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Sample/req
      -- CP-element group 34: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:next_ifetch_state_1358_936_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(34), ack => next_ifetch_state_1358_936_buf_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_update_start_
      -- CP-element group 35: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Update/req
      -- CP-element group 35: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:next_ifetch_state_1358_936_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(35), ack => next_ifetch_state_1358_936_buf_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Sample/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:next_ifetch_state_1358_936_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_ifetch_state_1358_936_buf_ack_0, ack => processor_daemon_CP_891_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_next_ifetch_state_936_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:next_ifetch_state_1358_936_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_ifetch_state_1358_936_buf_ack_1, ack => processor_daemon_CP_891_elements(37)); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	15 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(16);
      gj_processor_daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	13 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	200 
    -- CP-element group 39: 	172 
    -- CP-element group 39: 	176 
    -- CP-element group 39: 	208 
    -- CP-element group 39: 	160 
    -- CP-element group 39: 	168 
    -- CP-element group 39: 	152 
    -- CP-element group 39: 	156 
    -- CP-element group 39: 	184 
    -- CP-element group 39: 	188 
    -- CP-element group 39: 	192 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	17 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(200) & processor_daemon_CP_891_elements(172) & processor_daemon_CP_891_elements(176) & processor_daemon_CP_891_elements(208) & processor_daemon_CP_891_elements(160) & processor_daemon_CP_891_elements(168) & processor_daemon_CP_891_elements(152) & processor_daemon_CP_891_elements(156) & processor_daemon_CP_891_elements(184) & processor_daemon_CP_891_elements(188) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	15 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(40) <= processor_daemon_CP_891_elements(15);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	16 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	17 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(42) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(42) <= processor_daemon_CP_891_elements(17);
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	198 
    -- CP-element group 43: 	170 
    -- CP-element group 43: 	174 
    -- CP-element group 43: 	206 
    -- CP-element group 43: 	166 
    -- CP-element group 43: 	150 
    -- CP-element group 43: 	154 
    -- CP-element group 43: 	158 
    -- CP-element group 43: 	182 
    -- CP-element group 43: 	186 
    -- CP-element group 43: 	190 
    -- CP-element group 43: 	18 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	11 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_loopback_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(44) <= processor_daemon_CP_891_elements(11);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_loopback_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_937_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_937_loopback_sample_req_1041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_937_loopback_sample_req_1041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(45), ack => phi_stmt_937_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	12 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_entry_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(46) <= processor_daemon_CP_891_elements(12);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_entry_sample_req
      -- CP-element group 47: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_entry_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_937_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_937_entry_sample_req_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_937_entry_sample_req_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(47), ack => phi_stmt_937_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_phi_mux_ack_ps
      -- CP-element group 48: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_937_phi_mux_ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_937_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_937_phi_mux_ack_1047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_937_ack_0, ack => processor_daemon_CP_891_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_update_start_
      -- CP-element group 50: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(50) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(51) <= processor_daemon_CP_891_elements(52);
    -- CP-element group 52:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	51 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_939_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(52) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(52) is a control-delay.
    cp_element_52_delay: control_delay_element  generic map(name => " 52_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(50), ack => processor_daemon_CP_891_elements(52), clk => clk, reset =>reset);
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Sample/req
      -- CP-element group 53: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_icache_state_998_940_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(53), ack => n_icache_state_998_940_buf_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Update/req
      -- CP-element group 54: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_update_start_
      -- CP-element group 54: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_icache_state_998_940_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(54), ack => n_icache_state_998_940_buf_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_icache_state_998_940_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_icache_state_998_940_buf_ack_0, ack => processor_daemon_CP_891_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_icache_state_940_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_icache_state_998_940_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_icache_state_998_940_buf_ack_1, ack => processor_daemon_CP_891_elements(56)); -- 
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	161 
    -- CP-element group 57: 	165 
    -- CP-element group 57: 	169 
    -- CP-element group 57: 	153 
    -- CP-element group 57: 	157 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	15 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(57) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(161) & processor_daemon_CP_891_elements(165) & processor_daemon_CP_891_elements(169) & processor_daemon_CP_891_elements(153) & processor_daemon_CP_891_elements(157);
      gj_processor_daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	13 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	200 
    -- CP-element group 58: 	172 
    -- CP-element group 58: 	176 
    -- CP-element group 58: 	208 
    -- CP-element group 58: 	160 
    -- CP-element group 58: 	164 
    -- CP-element group 58: 	156 
    -- CP-element group 58: 	184 
    -- CP-element group 58: 	188 
    -- CP-element group 58: 	192 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	17 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(58) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(200) & processor_daemon_CP_891_elements(172) & processor_daemon_CP_891_elements(176) & processor_daemon_CP_891_elements(208) & processor_daemon_CP_891_elements(160) & processor_daemon_CP_891_elements(164) & processor_daemon_CP_891_elements(156) & processor_daemon_CP_891_elements(184) & processor_daemon_CP_891_elements(188) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	15 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(59) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(59) <= processor_daemon_CP_891_elements(15);
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(60) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	17 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(61) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(61) <= processor_daemon_CP_891_elements(17);
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	198 
    -- CP-element group 62: 	170 
    -- CP-element group 62: 	174 
    -- CP-element group 62: 	206 
    -- CP-element group 62: 	162 
    -- CP-element group 62: 	154 
    -- CP-element group 62: 	158 
    -- CP-element group 62: 	182 
    -- CP-element group 62: 	186 
    -- CP-element group 62: 	190 
    -- CP-element group 62: 	18 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_update_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(62) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	11 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_loopback_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(63) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(63) <= processor_daemon_CP_891_elements(11);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_loopback_sample_req_ps
      -- CP-element group 64: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_loopback_sample_req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_941_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_941_loopback_sample_req_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_941_loopback_sample_req_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(64), ack => phi_stmt_941_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_entry_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(65) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(65) <= processor_daemon_CP_891_elements(12);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_entry_sample_req_ps
      -- CP-element group 66: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_entry_sample_req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_941_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_941_entry_sample_req_1088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_941_entry_sample_req_1088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(66), ack => phi_stmt_941_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_phi_mux_ack_ps
      -- CP-element group 67: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_941_phi_mux_ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_941_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_941_phi_mux_ack_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_941_ack_0, ack => processor_daemon_CP_891_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(68) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_update_start_
      -- CP-element group 69: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(69) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(70) <= processor_daemon_CP_891_elements(71);
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	70 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_943_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(69), ack => processor_daemon_CP_891_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Sample/req
      -- CP-element group 72: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_idecode_state_1021_944_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(72), ack => n_idecode_state_1021_944_buf_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Update/req
      -- CP-element group 73: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_update_start_
      -- CP-element group 73: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_idecode_state_1021_944_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(73), ack => n_idecode_state_1021_944_buf_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Sample/ack
      -- CP-element group 74: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_idecode_state_1021_944_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_idecode_state_1021_944_buf_ack_0, ack => processor_daemon_CP_891_elements(74)); -- 
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Update/ack
      -- CP-element group 75: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_idecode_state_944_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_idecode_state_1021_944_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_idecode_state_1021_944_buf_ack_1, ack => processor_daemon_CP_891_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	13 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	16 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	15 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(76) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(16);
      gj_processor_daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	13 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	200 
    -- CP-element group 77: 	172 
    -- CP-element group 77: 	176 
    -- CP-element group 77: 	208 
    -- CP-element group 77: 	212 
    -- CP-element group 77: 	216 
    -- CP-element group 77: 	160 
    -- CP-element group 77: 	156 
    -- CP-element group 77: 	184 
    -- CP-element group 77: 	188 
    -- CP-element group 77: 	192 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	17 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(77) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(200) & processor_daemon_CP_891_elements(172) & processor_daemon_CP_891_elements(176) & processor_daemon_CP_891_elements(208) & processor_daemon_CP_891_elements(212) & processor_daemon_CP_891_elements(216) & processor_daemon_CP_891_elements(160) & processor_daemon_CP_891_elements(156) & processor_daemon_CP_891_elements(184) & processor_daemon_CP_891_elements(188) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	15 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(78) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(78) <= processor_daemon_CP_891_elements(15);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	16 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(79) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(80) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(80) <= processor_daemon_CP_891_elements(17);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	198 
    -- CP-element group 81: 	170 
    -- CP-element group 81: 	174 
    -- CP-element group 81: 	206 
    -- CP-element group 81: 	210 
    -- CP-element group 81: 	214 
    -- CP-element group 81: 	154 
    -- CP-element group 81: 	158 
    -- CP-element group 81: 	182 
    -- CP-element group 81: 	186 
    -- CP-element group 81: 	190 
    -- CP-element group 81: 	18 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(81) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	11 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_loopback_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(82) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(82) <= processor_daemon_CP_891_elements(11);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_loopback_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_945_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_945_loopback_sample_req_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_945_loopback_sample_req_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(83), ack => phi_stmt_945_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	12 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_entry_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(84) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(84) <= processor_daemon_CP_891_elements(12);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_entry_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_945_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_945_entry_sample_req_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_945_entry_sample_req_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(85), ack => phi_stmt_945_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_945_phi_mux_ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_945_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_945_phi_mux_ack_1135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_945_ack_0, ack => processor_daemon_CP_891_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(87) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(88) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(89) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(89) <= processor_daemon_CP_891_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_947_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(90) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(88), ack => processor_daemon_CP_891_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_sample_start__ps
      -- CP-element group 91: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iregfile_state_1030_948_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(91), ack => n_iregfile_state_1030_948_buf_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_update_start__ps
      -- CP-element group 92: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_update_start_
      -- CP-element group 92: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iregfile_state_1030_948_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(92), ack => n_iregfile_state_1030_948_buf_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_sample_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iregfile_state_1030_948_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iregfile_state_1030_948_buf_ack_0, ack => processor_daemon_CP_891_elements(93)); -- 
    -- CP-element group 94:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_update_completed__ps
      -- CP-element group 94: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iregfile_state_948_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iregfile_state_1030_948_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iregfile_state_1030_948_buf_ack_1, ack => processor_daemon_CP_891_elements(94)); -- 
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	13 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	16 
    -- CP-element group 95: 	193 
    -- CP-element group 95: 	197 
    -- CP-element group 95: 	201 
    -- CP-element group 95: 	205 
    -- CP-element group 95: 	209 
    -- CP-element group 95: 	213 
    -- CP-element group 95: 	217 
    -- CP-element group 95: 	189 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	15 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(95) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(193) & processor_daemon_CP_891_elements(197) & processor_daemon_CP_891_elements(201) & processor_daemon_CP_891_elements(205) & processor_daemon_CP_891_elements(209) & processor_daemon_CP_891_elements(213) & processor_daemon_CP_891_elements(217) & processor_daemon_CP_891_elements(189);
      gj_processor_daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	13 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	200 
    -- CP-element group 96: 	172 
    -- CP-element group 96: 	176 
    -- CP-element group 96: 	208 
    -- CP-element group 96: 	160 
    -- CP-element group 96: 	156 
    -- CP-element group 96: 	184 
    -- CP-element group 96: 	188 
    -- CP-element group 96: 	192 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	17 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(96) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 36) := "processor_daemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(200) & processor_daemon_CP_891_elements(172) & processor_daemon_CP_891_elements(176) & processor_daemon_CP_891_elements(208) & processor_daemon_CP_891_elements(160) & processor_daemon_CP_891_elements(156) & processor_daemon_CP_891_elements(184) & processor_daemon_CP_891_elements(188) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	15 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(97) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(97) <= processor_daemon_CP_891_elements(15);
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	16 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(98) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	17 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(99) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(99) <= processor_daemon_CP_891_elements(17);
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	198 
    -- CP-element group 100: 	170 
    -- CP-element group 100: 	174 
    -- CP-element group 100: 	206 
    -- CP-element group 100: 	154 
    -- CP-element group 100: 	158 
    -- CP-element group 100: 	182 
    -- CP-element group 100: 	186 
    -- CP-element group 100: 	190 
    -- CP-element group 100: 	18 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(100) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	11 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_loopback_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(101) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(101) <= processor_daemon_CP_891_elements(11);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_loopback_sample_req
      -- CP-element group 102: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_loopback_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_949_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_949_loopback_sample_req_1173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_949_loopback_sample_req_1173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(102), ack => phi_stmt_949_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	12 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_entry_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(103) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(103) <= processor_daemon_CP_891_elements(12);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_entry_sample_req
      -- CP-element group 104: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_entry_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_949_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_949_entry_sample_req_1176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_949_entry_sample_req_1176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(104), ack => phi_stmt_949_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_phi_mux_ack
      -- CP-element group 105: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_949_phi_mux_ack_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_949_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_949_phi_mux_ack_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_949_ack_0, ack => processor_daemon_CP_891_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(106) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(107) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(108) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(108) <= processor_daemon_CP_891_elements(109);
    -- CP-element group 109:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	108 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_951_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(109) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(107), ack => processor_daemon_CP_891_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_sample_start__ps
      -- CP-element group 110: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iexec_state_1275_952_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(110), ack => n_iexec_state_1275_952_buf_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_update_start__ps
      -- CP-element group 111: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_update_start_
      -- CP-element group 111: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iexec_state_1275_952_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(111), ack => n_iexec_state_1275_952_buf_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iexec_state_1275_952_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iexec_state_1275_952_buf_ack_0, ack => processor_daemon_CP_891_elements(112)); -- 
    -- CP-element group 113:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iexec_state_952_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iexec_state_1275_952_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iexec_state_1275_952_buf_ack_1, ack => processor_daemon_CP_891_elements(113)); -- 
    -- CP-element group 114:  join  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	13 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	16 
    -- CP-element group 114: 	181 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	15 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(114) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(181);
      gj_processor_daemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	13 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	200 
    -- CP-element group 115: 	172 
    -- CP-element group 115: 	176 
    -- CP-element group 115: 	228 
    -- CP-element group 115: 	232 
    -- CP-element group 115: 	236 
    -- CP-element group 115: 	208 
    -- CP-element group 115: 	220 
    -- CP-element group 115: 	224 
    -- CP-element group 115: 	160 
    -- CP-element group 115: 	156 
    -- CP-element group 115: 	184 
    -- CP-element group 115: 	188 
    -- CP-element group 115: 	192 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	17 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(115) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 14) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_markings: IntegerArray(0 to 14)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_delays: IntegerArray(0 to 14) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 15); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(200) & processor_daemon_CP_891_elements(172) & processor_daemon_CP_891_elements(176) & processor_daemon_CP_891_elements(228) & processor_daemon_CP_891_elements(232) & processor_daemon_CP_891_elements(236) & processor_daemon_CP_891_elements(208) & processor_daemon_CP_891_elements(220) & processor_daemon_CP_891_elements(224) & processor_daemon_CP_891_elements(160) & processor_daemon_CP_891_elements(156) & processor_daemon_CP_891_elements(184) & processor_daemon_CP_891_elements(188) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 15, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	15 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_sample_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(116) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(116) <= processor_daemon_CP_891_elements(15);
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	16 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(117) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	17 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_update_start__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(118) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(118) <= processor_daemon_CP_891_elements(17);
    -- CP-element group 119:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	198 
    -- CP-element group 119: 	170 
    -- CP-element group 119: 	174 
    -- CP-element group 119: 	230 
    -- CP-element group 119: 	234 
    -- CP-element group 119: 	206 
    -- CP-element group 119: 	218 
    -- CP-element group 119: 	222 
    -- CP-element group 119: 	226 
    -- CP-element group 119: 	154 
    -- CP-element group 119: 	158 
    -- CP-element group 119: 	182 
    -- CP-element group 119: 	186 
    -- CP-element group 119: 	190 
    -- CP-element group 119: 	18 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(119) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	11 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_loopback_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(120) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(120) <= processor_daemon_CP_891_elements(11);
    -- CP-element group 121:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_loopback_sample_req
      -- CP-element group 121: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_loopback_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_953_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_953_loopback_sample_req_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_953_loopback_sample_req_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(121), ack => phi_stmt_953_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	12 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_entry_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(122) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(122) <= processor_daemon_CP_891_elements(12);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_entry_sample_req
      -- CP-element group 123: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_entry_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_953_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_953_entry_sample_req_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_953_entry_sample_req_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(123), ack => phi_stmt_953_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_phi_mux_ack
      -- CP-element group 124: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_953_phi_mux_ack_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_953_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_953_phi_mux_ack_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_953_ack_0, ack => processor_daemon_CP_891_elements(124)); -- 
    -- CP-element group 125:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_sample_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(125) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(126) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(127) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(127) <= processor_daemon_CP_891_elements(128);
    -- CP-element group 128:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	127 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_955_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(128) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(128) is a control-delay.
    cp_element_128_delay: control_delay_element  generic map(name => " 128_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(126), ack => processor_daemon_CP_891_elements(128), clk => clk, reset =>reset);
    -- CP-element group 129:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (4) 
      -- CP-element group 129: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_sample_start__ps
      -- CP-element group 129: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_dcache_state_1142_956_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(129), ack => n_dcache_state_1142_956_buf_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (4) 
      -- CP-element group 130: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_update_start__ps
      -- CP-element group 130: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_update_start_
      -- CP-element group 130: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_dcache_state_1142_956_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(130), ack => n_dcache_state_1142_956_buf_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_sample_completed__ps
      -- CP-element group 131: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_dcache_state_1142_956_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_dcache_state_1142_956_buf_ack_0, ack => processor_daemon_CP_891_elements(131)); -- 
    -- CP-element group 132:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_update_completed__ps
      -- CP-element group 132: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_dcache_state_956_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_dcache_state_1142_956_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_dcache_state_1142_956_buf_ack_1, ack => processor_daemon_CP_891_elements(132)); -- 
    -- CP-element group 133:  join  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	16 
    -- CP-element group 133: 	229 
    -- CP-element group 133: 	233 
    -- CP-element group 133: 	237 
    -- CP-element group 133: 	221 
    -- CP-element group 133: 	225 
    -- CP-element group 133: 	185 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	15 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(133) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(229) & processor_daemon_CP_891_elements(233) & processor_daemon_CP_891_elements(237) & processor_daemon_CP_891_elements(221) & processor_daemon_CP_891_elements(225) & processor_daemon_CP_891_elements(185);
      gj_processor_daemon_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  join  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	13 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	239 
    -- CP-element group 134: 	196 
    -- CP-element group 134: 	200 
    -- CP-element group 134: 	172 
    -- CP-element group 134: 	176 
    -- CP-element group 134: 	204 
    -- CP-element group 134: 	208 
    -- CP-element group 134: 	160 
    -- CP-element group 134: 	156 
    -- CP-element group 134: 	184 
    -- CP-element group 134: 	188 
    -- CP-element group 134: 	192 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	17 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(134) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(13) & processor_daemon_CP_891_elements(239) & processor_daemon_CP_891_elements(196) & processor_daemon_CP_891_elements(200) & processor_daemon_CP_891_elements(172) & processor_daemon_CP_891_elements(176) & processor_daemon_CP_891_elements(204) & processor_daemon_CP_891_elements(208) & processor_daemon_CP_891_elements(160) & processor_daemon_CP_891_elements(156) & processor_daemon_CP_891_elements(184) & processor_daemon_CP_891_elements(188) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	16 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_sample_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(135) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(135) is bound as output of CP function.
    -- CP-element group 136:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	238 
    -- CP-element group 136: 	194 
    -- CP-element group 136: 	198 
    -- CP-element group 136: 	202 
    -- CP-element group 136: 	170 
    -- CP-element group 136: 	174 
    -- CP-element group 136: 	206 
    -- CP-element group 136: 	154 
    -- CP-element group 136: 	158 
    -- CP-element group 136: 	182 
    -- CP-element group 136: 	186 
    -- CP-element group 136: 	190 
    -- CP-element group 136: 	18 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(136) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_loopback_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(137) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(137) <= processor_daemon_CP_891_elements(11);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_loopback_sample_req
      -- CP-element group 138: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_loopback_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_957_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_957_loopback_sample_req_1261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_957_loopback_sample_req_1261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(138), ack => phi_stmt_957_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	12 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_entry_trigger
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(139) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(139) <= processor_daemon_CP_891_elements(12);
    -- CP-element group 140:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_entry_sample_req
      -- CP-element group 140: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_entry_sample_req_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_957_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_957_entry_sample_req_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_957_entry_sample_req_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(140), ack => phi_stmt_957_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_phi_mux_ack
      -- CP-element group 141: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/phi_stmt_957_phi_mux_ack_ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:phi_stmt_957_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_957_phi_mux_ack_1267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_957_ack_0, ack => processor_daemon_CP_891_elements(141)); -- 
    -- CP-element group 142:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_sample_start__ps
      -- CP-element group 142: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_sample_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(142) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(142) is bound as output of CP function.
    -- CP-element group 143:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_update_start__ps
      -- CP-element group 143: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(143) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(143) is bound as output of CP function.
    -- CP-element group 144:  join  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	145 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_update_completed__ps
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(144) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(144) <= processor_daemon_CP_891_elements(145);
    -- CP-element group 145:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	144 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/konst_959_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(145) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(145) is a control-delay.
    cp_element_145_delay: control_delay_element  generic map(name => " 145_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(143), ack => processor_daemon_CP_891_elements(145), clk => clk, reset =>reset);
    -- CP-element group 146:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iRetire_state_1317_960_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(146), ack => n_iRetire_state_1317_960_buf_req_0); -- 
    -- Element group processor_daemon_CP_891_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_update_start_
      -- CP-element group 147: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iRetire_state_1317_960_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(147), ack => n_iRetire_state_1317_960_buf_req_1); -- 
    -- Element group processor_daemon_CP_891_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (4) 
      -- CP-element group 148: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_sample_completed__ps
      -- CP-element group 148: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iRetire_state_1317_960_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iRetire_state_1317_960_buf_ack_0, ack => processor_daemon_CP_891_elements(148)); -- 
    -- CP-element group 149:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_update_completed__ps
      -- CP-element group 149: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/R_n_iRetire_state_960_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:n_iRetire_state_1317_960_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iRetire_state_1317_960_buf_ack_1, ack => processor_daemon_CP_891_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	43 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: 	185 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Sample/crr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_989_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(150), ack => call_stmt_989_call_req_0); -- 
    processor_daemon_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(152) & processor_daemon_CP_891_elements(185);
      gj_processor_daemon_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	16 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_update_start_
      -- CP-element group 151: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Update/ccr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_989_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(151), ack => call_stmt_989_call_req_1); -- 
    processor_daemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(153);
      gj_processor_daemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: 	39 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Sample/cra
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_989_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_989_call_ack_0, ack => processor_daemon_CP_891_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	242 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: 	57 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_Update/cca
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_989_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_989_call_ack_1, ack => processor_daemon_CP_891_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	136 
    -- CP-element group 154: 	119 
    -- CP-element group 154: 	24 
    -- CP-element group 154: 	43 
    -- CP-element group 154: 	62 
    -- CP-element group 154: 	81 
    -- CP-element group 154: 	100 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_idecode_1058_delayed_7_0_999_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(154), ack => W_flush_idecode_1058_delayed_7_0_999_inst_req_0); -- 
    processor_daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(156);
      gj_processor_daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	16 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_update_start_
      -- CP-element group 155: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_idecode_1058_delayed_7_0_999_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(155), ack => W_flush_idecode_1058_delayed_7_0_999_inst_req_1); -- 
    processor_daemon_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(157);
      gj_processor_daemon_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	134 
    -- CP-element group 156: 	115 
    -- CP-element group 156: 	154 
    -- CP-element group 156: 	20 
    -- CP-element group 156: 	39 
    -- CP-element group 156: 	58 
    -- CP-element group 156: 	77 
    -- CP-element group 156: 	96 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_idecode_1058_delayed_7_0_999_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_flush_idecode_1058_delayed_7_0_999_inst_ack_0, ack => processor_daemon_CP_891_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	243 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: 	57 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1001_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_idecode_1058_delayed_7_0_999_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_flush_idecode_1058_delayed_7_0_999_inst_ack_1, ack => processor_daemon_CP_891_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	136 
    -- CP-element group 158: 	119 
    -- CP-element group 158: 	24 
    -- CP-element group 158: 	43 
    -- CP-element group 158: 	62 
    -- CP-element group 158: 	81 
    -- CP-element group 158: 	100 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_stall_first_4_1060_delayed_7_0_1002_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(158), ack => W_stall_first_4_1060_delayed_7_0_1002_inst_req_0); -- 
    processor_daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(160);
      gj_processor_daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	16 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_update_start_
      -- CP-element group 159: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_stall_first_4_1060_delayed_7_0_1002_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(159), ack => W_stall_first_4_1060_delayed_7_0_1002_inst_req_1); -- 
    processor_daemon_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(161);
      gj_processor_daemon_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	134 
    -- CP-element group 160: 	115 
    -- CP-element group 160: 	158 
    -- CP-element group 160: 	20 
    -- CP-element group 160: 	39 
    -- CP-element group 160: 	58 
    -- CP-element group 160: 	77 
    -- CP-element group 160: 	96 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_stall_first_4_1060_delayed_7_0_1002_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_stall_first_4_1060_delayed_7_0_1002_inst_ack_0, ack => processor_daemon_CP_891_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	243 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	57 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1004_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_stall_first_4_1060_delayed_7_0_1002_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_stall_first_4_1060_delayed_7_0_1002_inst_ack_1, ack => processor_daemon_CP_891_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	62 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_idecode_state_1061_delayed_7_0_1005_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(162), ack => W_idecode_state_1061_delayed_7_0_1005_inst_req_0); -- 
    processor_daemon_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(164);
      gj_processor_daemon_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	16 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_update_start_
      -- CP-element group 163: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_idecode_state_1061_delayed_7_0_1005_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(163), ack => W_idecode_state_1061_delayed_7_0_1005_inst_req_1); -- 
    processor_daemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(165);
      gj_processor_daemon_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: 	58 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_idecode_state_1061_delayed_7_0_1005_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_idecode_state_1061_delayed_7_0_1005_inst_ack_0, ack => processor_daemon_CP_891_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	243 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	57 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1007_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_idecode_state_1061_delayed_7_0_1005_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_idecode_state_1061_delayed_7_0_1005_inst_ack_1, ack => processor_daemon_CP_891_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	43 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_icache_state_1063_delayed_7_0_1008_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(166), ack => W_icache_state_1063_delayed_7_0_1008_inst_req_0); -- 
    processor_daemon_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(168);
      gj_processor_daemon_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	16 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_update_start_
      -- CP-element group 167: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_icache_state_1063_delayed_7_0_1008_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(167), ack => W_icache_state_1063_delayed_7_0_1008_inst_req_1); -- 
    processor_daemon_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(169);
      gj_processor_daemon_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: 	39 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_icache_state_1063_delayed_7_0_1008_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_icache_state_1063_delayed_7_0_1008_inst_ack_0, ack => processor_daemon_CP_891_elements(168)); -- 
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	243 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	57 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1010_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_icache_state_1063_delayed_7_0_1008_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_icache_state_1063_delayed_7_0_1008_inst_ack_1, ack => processor_daemon_CP_891_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	136 
    -- CP-element group 170: 	119 
    -- CP-element group 170: 	24 
    -- CP-element group 170: 	43 
    -- CP-element group 170: 	62 
    -- CP-element group 170: 	81 
    -- CP-element group 170: 	100 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Sample/crr
      -- CP-element group 170: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Sample/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1133_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(170), ack => call_stmt_1133_call_req_0); -- 
    processor_daemon_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(172);
      gj_processor_daemon_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	180 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_update_start_
      -- CP-element group 171: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Update/ccr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1133_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(171), ack => call_stmt_1133_call_req_1); -- 
    processor_daemon_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= processor_daemon_CP_891_elements(180);
      gj_processor_daemon_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	134 
    -- CP-element group 172: 	170 
    -- CP-element group 172: 	115 
    -- CP-element group 172: 	20 
    -- CP-element group 172: 	39 
    -- CP-element group 172: 	58 
    -- CP-element group 172: 	77 
    -- CP-element group 172: 	96 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Sample/cra
      -- CP-element group 172: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Sample/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1133_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1133_call_ack_0, ack => processor_daemon_CP_891_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	178 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1133_Update/cca
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1133_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1133_call_ack_1, ack => processor_daemon_CP_891_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	136 
    -- CP-element group 174: 	119 
    -- CP-element group 174: 	24 
    -- CP-element group 174: 	43 
    -- CP-element group 174: 	62 
    -- CP-element group 174: 	81 
    -- CP-element group 174: 	100 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Sample/req
      -- CP-element group 174: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_dcache_1221_delayed_4_0_1134_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(174), ack => W_flush_dcache_1221_delayed_4_0_1134_inst_req_0); -- 
    processor_daemon_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(176);
      gj_processor_daemon_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	180 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_update_start_
      -- CP-element group 175: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Update/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_dcache_1221_delayed_4_0_1134_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(175), ack => W_flush_dcache_1221_delayed_4_0_1134_inst_req_1); -- 
    processor_daemon_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= processor_daemon_CP_891_elements(180);
      gj_processor_daemon_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	134 
    -- CP-element group 176: 	174 
    -- CP-element group 176: 	115 
    -- CP-element group 176: 	20 
    -- CP-element group 176: 	39 
    -- CP-element group 176: 	58 
    -- CP-element group 176: 	77 
    -- CP-element group 176: 	96 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_dcache_1221_delayed_4_0_1134_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_flush_dcache_1221_delayed_4_0_1134_inst_ack_0, ack => processor_daemon_CP_891_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1136_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_dcache_1221_delayed_4_0_1134_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_flush_dcache_1221_delayed_4_0_1134_inst_ack_1, ack => processor_daemon_CP_891_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	173 
    -- CP-element group 178: 	177 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_start/$entry
      -- CP-element group 178: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_start/req
      -- CP-element group 178: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:MUX_1141_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(178), ack => MUX_1141_inst_req_0); -- 
    processor_daemon_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(173) & processor_daemon_CP_891_elements(177) & processor_daemon_CP_891_elements(180);
      gj_processor_daemon_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	16 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_complete/req
      -- CP-element group 179: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_update_start_
      -- CP-element group 179: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_complete/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:MUX_1141_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(179), ack => MUX_1141_inst_req_1); -- 
    processor_daemon_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(181);
      gj_processor_daemon_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	171 
    -- CP-element group 180: 	175 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_start/ack
      -- CP-element group 180: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_start/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:MUX_1141_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1141_inst_ack_0, ack => processor_daemon_CP_891_elements(180)); -- 
    -- CP-element group 181:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	243 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: 	114 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_complete/ack
      -- CP-element group 181: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/MUX_1141_complete/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:MUX_1141_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1141_inst_ack_1, ack => processor_daemon_CP_891_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	136 
    -- CP-element group 182: 	242 
    -- CP-element group 182: 	119 
    -- CP-element group 182: 	24 
    -- CP-element group 182: 	43 
    -- CP-element group 182: 	62 
    -- CP-element group 182: 	81 
    -- CP-element group 182: 	100 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Sample/crr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1175_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(182), ack => call_stmt_1175_call_req_0); -- 
    processor_daemon_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(242) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(184);
      gj_processor_daemon_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	16 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_update_start_
      -- CP-element group 183: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Update/ccr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1175_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(183), ack => call_stmt_1175_call_req_1); -- 
    processor_daemon_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(185);
      gj_processor_daemon_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	134 
    -- CP-element group 184: 	115 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	20 
    -- CP-element group 184: 	39 
    -- CP-element group 184: 	58 
    -- CP-element group 184: 	77 
    -- CP-element group 184: 	96 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Sample/cra
      -- CP-element group 184: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Sample/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1175_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1175_call_ack_0, ack => processor_daemon_CP_891_elements(184)); -- 
    -- CP-element group 185:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	243 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	133 
    -- CP-element group 185: 	150 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (4) 
      -- CP-element group 185: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1175_Update/cca
      -- CP-element group 185: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/ring_reenable_memory_space_0
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1175_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1175_call_ack_1, ack => processor_daemon_CP_891_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	136 
    -- CP-element group 186: 	119 
    -- CP-element group 186: 	24 
    -- CP-element group 186: 	43 
    -- CP-element group 186: 	62 
    -- CP-element group 186: 	81 
    -- CP-element group 186: 	100 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Sample/crr
      -- CP-element group 186: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Sample/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(186) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1224_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(186), ack => call_stmt_1224_call_req_0); -- 
    processor_daemon_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(188);
      gj_processor_daemon_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	16 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	189 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_update_start_
      -- CP-element group 187: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Update/ccr
      -- CP-element group 187: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Update/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1224_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(187), ack => call_stmt_1224_call_req_1); -- 
    processor_daemon_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(189);
      gj_processor_daemon_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	134 
    -- CP-element group 188: 	115 
    -- CP-element group 188: 	186 
    -- CP-element group 188: 	20 
    -- CP-element group 188: 	39 
    -- CP-element group 188: 	58 
    -- CP-element group 188: 	77 
    -- CP-element group 188: 	96 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Sample/cra
      -- CP-element group 188: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Sample/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1224_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1224_call_ack_0, ack => processor_daemon_CP_891_elements(188)); -- 
    -- CP-element group 189:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	243 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: 	95 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Update/cca
      -- CP-element group 189: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_1224_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:call_stmt_1224_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1224_call_ack_1, ack => processor_daemon_CP_891_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	136 
    -- CP-element group 190: 	119 
    -- CP-element group 190: 	24 
    -- CP-element group 190: 	43 
    -- CP-element group 190: 	62 
    -- CP-element group 190: 	81 
    -- CP-element group 190: 	100 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Sample/req
      -- CP-element group 190: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(190), ack => W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_0); -- 
    processor_daemon_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(192);
      gj_processor_daemon_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	16 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Update/req
      -- CP-element group 191: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(191), ack => W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_1); -- 
    processor_daemon_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(193);
      gj_processor_daemon_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	134 
    -- CP-element group 192: 	115 
    -- CP-element group 192: 	190 
    -- CP-element group 192: 	20 
    -- CP-element group 192: 	39 
    -- CP-element group 192: 	58 
    -- CP-element group 192: 	77 
    -- CP-element group 192: 	96 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Sample/ack
      -- CP-element group 192: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(192) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_0, ack => processor_daemon_CP_891_elements(192)); -- 
    -- CP-element group 193:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	243 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: 	95 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_Update/ack
      -- CP-element group 193: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1227_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_1, ack => processor_daemon_CP_891_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	136 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Sample/req
      -- CP-element group 194: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(194), ack => W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_0); -- 
    processor_daemon_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(196);
      gj_processor_daemon_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	16 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	197 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Update/req
      -- CP-element group 195: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(195), ack => W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_1); -- 
    processor_daemon_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(197);
      gj_processor_daemon_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	134 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(196) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_0, ack => processor_daemon_CP_891_elements(196)); -- 
    -- CP-element group 197:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	243 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: 	95 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1230_Update/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(197)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(197)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(197) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_1, ack => processor_daemon_CP_891_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	136 
    -- CP-element group 198: 	119 
    -- CP-element group 198: 	24 
    -- CP-element group 198: 	43 
    -- CP-element group 198: 	62 
    -- CP-element group 198: 	81 
    -- CP-element group 198: 	100 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Sample/req
      -- CP-element group 198: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(198)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(198)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(198) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(198), ack => W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_0); -- 
    processor_daemon_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(200);
      gj_processor_daemon_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	16 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	201 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Update/req
      -- CP-element group 199: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_update_start_
      -- CP-element group 199: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Update/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(199)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(199)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(199) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(199), ack => W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_1); -- 
    processor_daemon_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(201);
      gj_processor_daemon_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	134 
    -- CP-element group 200: 	198 
    -- CP-element group 200: 	115 
    -- CP-element group 200: 	20 
    -- CP-element group 200: 	39 
    -- CP-element group 200: 	58 
    -- CP-element group 200: 	77 
    -- CP-element group 200: 	96 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Sample/ack
      -- CP-element group 200: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(200)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(200)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(200) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_0, ack => processor_daemon_CP_891_elements(200)); -- 
    -- CP-element group 201:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	243 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: 	95 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Update/ack
      -- CP-element group 201: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1239_Update/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(201)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(201)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(201) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_1, ack => processor_daemon_CP_891_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	136 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Sample/req
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(202)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(202)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(202) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(202), ack => W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_0); -- 
    processor_daemon_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(204);
      gj_processor_daemon_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	16 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_update_start_
      -- CP-element group 203: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Update/req
      -- CP-element group 203: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Update/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(203)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(203)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(203) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(203), ack => W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_1); -- 
    processor_daemon_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(205);
      gj_processor_daemon_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	134 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Sample/ack
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(204)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(204)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(204) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_0, ack => processor_daemon_CP_891_elements(204)); -- 
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	243 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: 	95 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Update/ack
      -- CP-element group 205: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1242_Update/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(205)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(205)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(205) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_1, ack => processor_daemon_CP_891_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	136 
    -- CP-element group 206: 	119 
    -- CP-element group 206: 	24 
    -- CP-element group 206: 	43 
    -- CP-element group 206: 	62 
    -- CP-element group 206: 	81 
    -- CP-element group 206: 	100 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Sample/req
      -- CP-element group 206: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Sample/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(206)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(206)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(206) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_iexec_1330_delayed_7_0_1249_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(206), ack => W_flush_iexec_1330_delayed_7_0_1249_inst_req_0); -- 
    processor_daemon_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(24) & processor_daemon_CP_891_elements(43) & processor_daemon_CP_891_elements(62) & processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(100) & processor_daemon_CP_891_elements(208);
      gj_processor_daemon_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	16 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_update_start_
      -- CP-element group 207: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Update/req
      -- CP-element group 207: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Update/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(207)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(207)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(207) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_iexec_1330_delayed_7_0_1249_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(207), ack => W_flush_iexec_1330_delayed_7_0_1249_inst_req_1); -- 
    processor_daemon_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(209);
      gj_processor_daemon_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	134 
    -- CP-element group 208: 	206 
    -- CP-element group 208: 	115 
    -- CP-element group 208: 	20 
    -- CP-element group 208: 	39 
    -- CP-element group 208: 	58 
    -- CP-element group 208: 	77 
    -- CP-element group 208: 	96 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Sample/ack
      -- CP-element group 208: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Sample/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(208)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(208)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(208) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_iexec_1330_delayed_7_0_1249_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_flush_iexec_1330_delayed_7_0_1249_inst_ack_0, ack => processor_daemon_CP_891_elements(208)); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	243 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: 	95 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Update/ack
      -- CP-element group 209: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1251_Update/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(209)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(209)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(209) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_flush_iexec_1330_delayed_7_0_1249_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_flush_iexec_1330_delayed_7_0_1249_inst_ack_1, ack => processor_daemon_CP_891_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	81 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Sample/rr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(210)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(210)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(210) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u16_u32_1259_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(210), ack => CONCAT_u16_u32_1259_inst_req_0); -- 
    processor_daemon_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(212);
      gj_processor_daemon_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	16 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_update_start_
      -- CP-element group 211: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Update/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(211)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(211)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(211) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u16_u32_1259_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(211), ack => CONCAT_u16_u32_1259_inst_req_1); -- 
    processor_daemon_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(213);
      gj_processor_daemon_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: 	77 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Sample/ra
      -- CP-element group 212: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(212)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(212)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(212) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u16_u32_1259_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1259_inst_ack_0, ack => processor_daemon_CP_891_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	243 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: 	95 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u16_u32_1259_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(213)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(213)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(213) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u16_u32_1259_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1259_inst_ack_1, ack => processor_daemon_CP_891_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	81 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Sample/req
      -- CP-element group 214: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Sample/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(214)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(214)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(214) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iregfile_pc_1342_delayed_7_0_1261_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(214), ack => W_iregfile_pc_1342_delayed_7_0_1261_inst_req_0); -- 
    processor_daemon_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(81) & processor_daemon_CP_891_elements(216);
      gj_processor_daemon_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	16 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	217 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_update_start_
      -- CP-element group 215: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Update/req
      -- CP-element group 215: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Update/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(215)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(215)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(215) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iregfile_pc_1342_delayed_7_0_1261_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(215), ack => W_iregfile_pc_1342_delayed_7_0_1261_inst_req_1); -- 
    processor_daemon_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(217);
      gj_processor_daemon_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: 	77 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Sample/ack
      -- CP-element group 216: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(216)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(216)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(216) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_0, ack => processor_daemon_CP_891_elements(216)); -- 
    -- CP-element group 217:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	243 
    -- CP-element group 217: marked-successors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: 	95 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Update/ack
      -- CP-element group 217: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1263_Update/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(217)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(217)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(217) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_1, ack => processor_daemon_CP_891_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	119 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(218)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(218)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(218) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:EQ_u8_u1_1279_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(218), ack => EQ_u8_u1_1279_inst_req_0); -- 
    processor_daemon_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(220);
      gj_processor_daemon_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	16 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Update/cr
      -- CP-element group 219: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(219)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(219)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(219) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:EQ_u8_u1_1279_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(219), ack => EQ_u8_u1_1279_inst_req_1); -- 
    processor_daemon_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(221);
      gj_processor_daemon_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: 	115 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Sample/ra
      -- CP-element group 220: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(220)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(220)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(220) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:EQ_u8_u1_1279_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_1279_inst_ack_0, ack => processor_daemon_CP_891_elements(220)); -- 
    -- CP-element group 221:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	243 
    -- CP-element group 221: marked-successors 
    -- CP-element group 221: 	133 
    -- CP-element group 221: 	219 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/EQ_u8_u1_1279_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(221)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(221)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(221) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:EQ_u8_u1_1279_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_1279_inst_ack_1, ack => processor_daemon_CP_891_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	119 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Sample/req
      -- CP-element group 222: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(222)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(222)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(222) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(222), ack => W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_0); -- 
    processor_daemon_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(224);
      gj_processor_daemon_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	16 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	225 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Update/req
      -- CP-element group 223: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(223)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(223)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(223) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(223), ack => W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_1); -- 
    processor_daemon_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(225);
      gj_processor_daemon_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: 	115 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Sample/ack
      -- CP-element group 224: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(224)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(224)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(224) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_0, ack => processor_daemon_CP_891_elements(224)); -- 
    -- CP-element group 225:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	243 
    -- CP-element group 225: marked-successors 
    -- CP-element group 225: 	133 
    -- CP-element group 225: 	223 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Update/ack
      -- CP-element group 225: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1283_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(225)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(225)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(225) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_1, ack => processor_daemon_CP_891_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	119 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Sample/rr
      -- CP-element group 226: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(226)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(226)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(226) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u24_u64_1299_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(226), ack => CONCAT_u24_u64_1299_inst_req_0); -- 
    processor_daemon_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(228);
      gj_processor_daemon_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	16 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	229 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_update_start_
      -- CP-element group 227: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Update/cr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(227)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(227)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(227) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u24_u64_1299_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(227), ack => CONCAT_u24_u64_1299_inst_req_1); -- 
    processor_daemon_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(229);
      gj_processor_daemon_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: 	115 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Sample/ra
      -- CP-element group 228: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(228)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(228)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(228) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u24_u64_1299_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u24_u64_1299_inst_ack_0, ack => processor_daemon_CP_891_elements(228)); -- 
    -- CP-element group 229:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	243 
    -- CP-element group 229: marked-successors 
    -- CP-element group 229: 	133 
    -- CP-element group 229: 	227 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Update/ca
      -- CP-element group 229: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u24_u64_1299_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(229)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(229)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(229) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u24_u64_1299_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u24_u64_1299_inst_ack_1, ack => processor_daemon_CP_891_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	119 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Sample/req
      -- CP-element group 230: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Sample/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(230)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(230)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(230) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_rd2_1365_delayed_7_0_1301_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(230), ack => W_dcache_rd2_1365_delayed_7_0_1301_inst_req_0); -- 
    processor_daemon_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(232);
      gj_processor_daemon_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	16 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	233 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	233 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Update/req
      -- CP-element group 231: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(231)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(231)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(231) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_rd2_1365_delayed_7_0_1301_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(231), ack => W_dcache_rd2_1365_delayed_7_0_1301_inst_req_1); -- 
    processor_daemon_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(233);
      gj_processor_daemon_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: 	115 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Sample/ack
      -- CP-element group 232: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(232)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(232)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(232) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_0, ack => processor_daemon_CP_891_elements(232)); -- 
    -- CP-element group 233:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	243 
    -- CP-element group 233: marked-successors 
    -- CP-element group 233: 	133 
    -- CP-element group 233: 	231 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Update/ack
      -- CP-element group 233: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/assign_stmt_1303_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(233)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(233)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(233) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_1, ack => processor_daemon_CP_891_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	119 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_sample_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(234)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(234)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(234) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u1_u11_1307_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(234), ack => CONCAT_u1_u11_1307_inst_req_0); -- 
    processor_daemon_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(119) & processor_daemon_CP_891_elements(236);
      gj_processor_daemon_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	16 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	237 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_update_start_
      -- CP-element group 235: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Update/cr
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(235)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(235)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(235) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u1_u11_1307_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(235), ack => CONCAT_u1_u11_1307_inst_req_1); -- 
    processor_daemon_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(237);
      gj_processor_daemon_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	115 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Sample/ra
      -- CP-element group 236: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_sample_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(236)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(236)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(236) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u1_u11_1307_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u11_1307_inst_ack_0, ack => processor_daemon_CP_891_elements(236)); -- 
    -- CP-element group 237:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	243 
    -- CP-element group 237: marked-successors 
    -- CP-element group 237: 	133 
    -- CP-element group 237: 	235 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_Update/ca
      -- CP-element group 237: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/CONCAT_u1_u11_1307_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(237)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(237)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(237) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:CONCAT_u1_u11_1307_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u11_1307_inst_ack_1, ack => processor_daemon_CP_891_elements(237)); -- 
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	136 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Sample/$entry
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(238)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(238)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(238) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:WPIPE_processor_result_1370_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(238), ack => WPIPE_processor_result_1370_inst_req_0); -- 
    processor_daemon_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(136) & processor_daemon_CP_891_elements(240);
      gj_processor_daemon_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	134 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Update/req
      -- CP-element group 239: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_update_start_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(239)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(239)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(239) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:WPIPE_processor_result_1370_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:WPIPE_processor_result_1370_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_processor_result_1370_inst_ack_0, ack => processor_daemon_CP_891_elements(239)); -- 
    req_1616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(239), ack => WPIPE_processor_result_1370_inst_req_1); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	243 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/WPIPE_processor_result_1370_update_completed_
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(240)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(240)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(240) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:WPIPE_processor_result_1370_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_processor_result_1370_inst_ack_1, ack => processor_daemon_CP_891_elements(240)); -- 
    -- CP-element group 241:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	13 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	14 
    -- CP-element group 241:  members (1) 
      -- CP-element group 241: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(241)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(241)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(241) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(241) is a control-delay.
    cp_element_241_delay: control_delay_element  generic map(name => " 241_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(13), ack => processor_daemon_CP_891_elements(241), clk => clk, reset =>reset);
    -- CP-element group 242:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	153 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	182 
    -- CP-element group 242:  members (1) 
      -- CP-element group 242: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/call_stmt_989_call_stmt_1175_delay
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(242)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(242)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(242) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processor_daemon_CP_891_elements(242) is a control-delay.
    cp_element_242_delay: control_delay_element  generic map(name => " 242_delay", delay_value => 1)  port map(req => processor_daemon_CP_891_elements(153), ack => processor_daemon_CP_891_elements(242), clk => clk, reset =>reset);
    -- CP-element group 243:  join  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	16 
    -- CP-element group 243: 	240 
    -- CP-element group 243: 	193 
    -- CP-element group 243: 	197 
    -- CP-element group 243: 	201 
    -- CP-element group 243: 	229 
    -- CP-element group 243: 	233 
    -- CP-element group 243: 	237 
    -- CP-element group 243: 	205 
    -- CP-element group 243: 	209 
    -- CP-element group 243: 	213 
    -- CP-element group 243: 	217 
    -- CP-element group 243: 	221 
    -- CP-element group 243: 	225 
    -- CP-element group 243: 	161 
    -- CP-element group 243: 	165 
    -- CP-element group 243: 	169 
    -- CP-element group 243: 	157 
    -- CP-element group 243: 	181 
    -- CP-element group 243: 	185 
    -- CP-element group 243: 	189 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	10 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/do_while_stmt_931_loop_body/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(243)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(243)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(243) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant joinName: string(1 to 37) := "processor_daemon_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= processor_daemon_CP_891_elements(16) & processor_daemon_CP_891_elements(240) & processor_daemon_CP_891_elements(193) & processor_daemon_CP_891_elements(197) & processor_daemon_CP_891_elements(201) & processor_daemon_CP_891_elements(229) & processor_daemon_CP_891_elements(233) & processor_daemon_CP_891_elements(237) & processor_daemon_CP_891_elements(205) & processor_daemon_CP_891_elements(209) & processor_daemon_CP_891_elements(213) & processor_daemon_CP_891_elements(217) & processor_daemon_CP_891_elements(221) & processor_daemon_CP_891_elements(225) & processor_daemon_CP_891_elements(161) & processor_daemon_CP_891_elements(165) & processor_daemon_CP_891_elements(169) & processor_daemon_CP_891_elements(157) & processor_daemon_CP_891_elements(181) & processor_daemon_CP_891_elements(185) & processor_daemon_CP_891_elements(189);
      gj_processor_daemon_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processor_daemon_CP_891_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	9 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (2) 
      -- CP-element group 244: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_exit/ack
      -- CP-element group 244: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_exit/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(244)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(244)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(244) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:do_while_stmt_931_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_931_branch_ack_0, ack => processor_daemon_CP_891_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	9 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (2) 
      -- CP-element group 245: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_taken/ack
      -- CP-element group 245: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/loop_taken/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(245)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(245)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(245) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:do_while_stmt_931_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_931_branch_ack_1, ack => processor_daemon_CP_891_elements(245)); -- 
    -- CP-element group 246:  transition  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	7 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	5 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_921/branch_block_stmt_930/do_while_stmt_931/$exit
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(246)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(246)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(246) fired."); 
        -- 
      end if; --
    end process; 
    processor_daemon_CP_891_elements(246) <= processor_daemon_CP_891_elements(7);
    -- CP-element group 247:  merge  transition  place  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	5 
    -- CP-element group 247: 	0 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	1 
    -- CP-element group 247:  members (10) 
      -- CP-element group 247: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_921/assign_stmt_925__entry__
      -- CP-element group 247: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_921/assign_stmt_925/$entry
      -- CP-element group 247: 	 branch_block_stmt_921/merge_stmt_922__exit__
      -- CP-element group 247: 	 branch_block_stmt_921/assign_stmt_925/RPIPE_start_processor_924_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_921/merge_stmt_922_PhiReqMerge
      -- CP-element group 247: 	 branch_block_stmt_921/merge_stmt_922_PhiAck/$entry
      -- CP-element group 247: 	 branch_block_stmt_921/merge_stmt_922_PhiAck/$exit
      -- CP-element group 247: 	 branch_block_stmt_921/merge_stmt_922_PhiAck/dummy
      -- 
    -- logger for CP element group processor_daemon_CP_891_elements(247)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processor_daemon_CP_891_elements(247)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:processor_daemon_CP_891_elements(247) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processor_daemon:CP:RPIPE_start_processor_924_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processor_daemon_CP_891_elements(247), ack => RPIPE_start_processor_924_inst_req_0); -- 
    processor_daemon_CP_891_elements(247) <= OrReduce(processor_daemon_CP_891_elements(5) & processor_daemon_CP_891_elements(0));
    processor_daemon_do_while_stmt_931_terminator_1629: loop_terminator -- 
      generic map (name => " processor_daemon_do_while_stmt_931_terminator_1629", max_iterations_in_flight =>15) 
      port map(loop_body_exit => processor_daemon_CP_891_elements(10),loop_continue => processor_daemon_CP_891_elements(245),loop_terminate => processor_daemon_CP_891_elements(244),loop_back => processor_daemon_CP_891_elements(8),loop_exit => processor_daemon_CP_891_elements(7),clk => clk, reset => reset); -- 
    phi_stmt_933_phi_seq_1031_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= processor_daemon_CP_891_elements(27);
      processor_daemon_CP_891_elements(30)<= src_sample_reqs(0);
      src_sample_acks(0)  <= processor_daemon_CP_891_elements(30);
      processor_daemon_CP_891_elements(31)<= src_update_reqs(0);
      src_update_acks(0)  <= processor_daemon_CP_891_elements(32);
      processor_daemon_CP_891_elements(28) <= phi_mux_reqs(0);
      triggers(1)  <= processor_daemon_CP_891_elements(25);
      processor_daemon_CP_891_elements(34)<= src_sample_reqs(1);
      src_sample_acks(1)  <= processor_daemon_CP_891_elements(36);
      processor_daemon_CP_891_elements(35)<= src_update_reqs(1);
      src_update_acks(1)  <= processor_daemon_CP_891_elements(37);
      processor_daemon_CP_891_elements(26) <= phi_mux_reqs(1);
      phi_stmt_933_phi_seq_1031 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_933_phi_seq_1031") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => processor_daemon_CP_891_elements(21), 
          phi_sample_ack => processor_daemon_CP_891_elements(22), 
          phi_update_req => processor_daemon_CP_891_elements(23), 
          phi_update_ack => processor_daemon_CP_891_elements(24), 
          phi_mux_ack => processor_daemon_CP_891_elements(29), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_937_phi_seq_1075_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= processor_daemon_CP_891_elements(46);
      processor_daemon_CP_891_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= processor_daemon_CP_891_elements(49);
      processor_daemon_CP_891_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= processor_daemon_CP_891_elements(51);
      processor_daemon_CP_891_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= processor_daemon_CP_891_elements(44);
      processor_daemon_CP_891_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= processor_daemon_CP_891_elements(55);
      processor_daemon_CP_891_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= processor_daemon_CP_891_elements(56);
      processor_daemon_CP_891_elements(45) <= phi_mux_reqs(1);
      phi_stmt_937_phi_seq_1075 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_937_phi_seq_1075") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => processor_daemon_CP_891_elements(40), 
          phi_sample_ack => processor_daemon_CP_891_elements(41), 
          phi_update_req => processor_daemon_CP_891_elements(42), 
          phi_update_ack => processor_daemon_CP_891_elements(43), 
          phi_mux_ack => processor_daemon_CP_891_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_941_phi_seq_1119_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= processor_daemon_CP_891_elements(65);
      processor_daemon_CP_891_elements(68)<= src_sample_reqs(0);
      src_sample_acks(0)  <= processor_daemon_CP_891_elements(68);
      processor_daemon_CP_891_elements(69)<= src_update_reqs(0);
      src_update_acks(0)  <= processor_daemon_CP_891_elements(70);
      processor_daemon_CP_891_elements(66) <= phi_mux_reqs(0);
      triggers(1)  <= processor_daemon_CP_891_elements(63);
      processor_daemon_CP_891_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= processor_daemon_CP_891_elements(74);
      processor_daemon_CP_891_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= processor_daemon_CP_891_elements(75);
      processor_daemon_CP_891_elements(64) <= phi_mux_reqs(1);
      phi_stmt_941_phi_seq_1119 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_941_phi_seq_1119") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => processor_daemon_CP_891_elements(59), 
          phi_sample_ack => processor_daemon_CP_891_elements(60), 
          phi_update_req => processor_daemon_CP_891_elements(61), 
          phi_update_ack => processor_daemon_CP_891_elements(62), 
          phi_mux_ack => processor_daemon_CP_891_elements(67), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_945_phi_seq_1163_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= processor_daemon_CP_891_elements(84);
      processor_daemon_CP_891_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= processor_daemon_CP_891_elements(87);
      processor_daemon_CP_891_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= processor_daemon_CP_891_elements(89);
      processor_daemon_CP_891_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= processor_daemon_CP_891_elements(82);
      processor_daemon_CP_891_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= processor_daemon_CP_891_elements(93);
      processor_daemon_CP_891_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= processor_daemon_CP_891_elements(94);
      processor_daemon_CP_891_elements(83) <= phi_mux_reqs(1);
      phi_stmt_945_phi_seq_1163 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_945_phi_seq_1163") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => processor_daemon_CP_891_elements(78), 
          phi_sample_ack => processor_daemon_CP_891_elements(79), 
          phi_update_req => processor_daemon_CP_891_elements(80), 
          phi_update_ack => processor_daemon_CP_891_elements(81), 
          phi_mux_ack => processor_daemon_CP_891_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_949_phi_seq_1207_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= processor_daemon_CP_891_elements(103);
      processor_daemon_CP_891_elements(106)<= src_sample_reqs(0);
      src_sample_acks(0)  <= processor_daemon_CP_891_elements(106);
      processor_daemon_CP_891_elements(107)<= src_update_reqs(0);
      src_update_acks(0)  <= processor_daemon_CP_891_elements(108);
      processor_daemon_CP_891_elements(104) <= phi_mux_reqs(0);
      triggers(1)  <= processor_daemon_CP_891_elements(101);
      processor_daemon_CP_891_elements(110)<= src_sample_reqs(1);
      src_sample_acks(1)  <= processor_daemon_CP_891_elements(112);
      processor_daemon_CP_891_elements(111)<= src_update_reqs(1);
      src_update_acks(1)  <= processor_daemon_CP_891_elements(113);
      processor_daemon_CP_891_elements(102) <= phi_mux_reqs(1);
      phi_stmt_949_phi_seq_1207 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_949_phi_seq_1207") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => processor_daemon_CP_891_elements(97), 
          phi_sample_ack => processor_daemon_CP_891_elements(98), 
          phi_update_req => processor_daemon_CP_891_elements(99), 
          phi_update_ack => processor_daemon_CP_891_elements(100), 
          phi_mux_ack => processor_daemon_CP_891_elements(105), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_953_phi_seq_1251_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= processor_daemon_CP_891_elements(122);
      processor_daemon_CP_891_elements(125)<= src_sample_reqs(0);
      src_sample_acks(0)  <= processor_daemon_CP_891_elements(125);
      processor_daemon_CP_891_elements(126)<= src_update_reqs(0);
      src_update_acks(0)  <= processor_daemon_CP_891_elements(127);
      processor_daemon_CP_891_elements(123) <= phi_mux_reqs(0);
      triggers(1)  <= processor_daemon_CP_891_elements(120);
      processor_daemon_CP_891_elements(129)<= src_sample_reqs(1);
      src_sample_acks(1)  <= processor_daemon_CP_891_elements(131);
      processor_daemon_CP_891_elements(130)<= src_update_reqs(1);
      src_update_acks(1)  <= processor_daemon_CP_891_elements(132);
      processor_daemon_CP_891_elements(121) <= phi_mux_reqs(1);
      phi_stmt_953_phi_seq_1251 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_953_phi_seq_1251") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => processor_daemon_CP_891_elements(116), 
          phi_sample_ack => processor_daemon_CP_891_elements(117), 
          phi_update_req => processor_daemon_CP_891_elements(118), 
          phi_update_ack => processor_daemon_CP_891_elements(119), 
          phi_mux_ack => processor_daemon_CP_891_elements(124), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_957_phi_seq_1295_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= processor_daemon_CP_891_elements(139);
      processor_daemon_CP_891_elements(142)<= src_sample_reqs(0);
      src_sample_acks(0)  <= processor_daemon_CP_891_elements(142);
      processor_daemon_CP_891_elements(143)<= src_update_reqs(0);
      src_update_acks(0)  <= processor_daemon_CP_891_elements(144);
      processor_daemon_CP_891_elements(140) <= phi_mux_reqs(0);
      triggers(1)  <= processor_daemon_CP_891_elements(137);
      processor_daemon_CP_891_elements(146)<= src_sample_reqs(1);
      src_sample_acks(1)  <= processor_daemon_CP_891_elements(148);
      processor_daemon_CP_891_elements(147)<= src_update_reqs(1);
      src_update_acks(1)  <= processor_daemon_CP_891_elements(149);
      processor_daemon_CP_891_elements(138) <= phi_mux_reqs(1);
      phi_stmt_957_phi_seq_1295 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_957_phi_seq_1295") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => processor_daemon_CP_891_elements(15), 
          phi_sample_ack => processor_daemon_CP_891_elements(135), 
          phi_update_req => processor_daemon_CP_891_elements(17), 
          phi_update_ack => processor_daemon_CP_891_elements(136), 
          phi_mux_ack => processor_daemon_CP_891_elements(141), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_983_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= processor_daemon_CP_891_elements(11);
        preds(1)  <= processor_daemon_CP_891_elements(12);
        entry_tmerge_983 : transition_merge -- 
          generic map(name => " entry_tmerge_983")
          port map (preds => preds, symbol_out => processor_daemon_CP_891_elements(13));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u10_u10_1349_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u16_u24_1295_wire : std_logic_vector(23 downto 0);
    signal CONCAT_u16_u32_1338_1338_delayed_7_0_1260 : std_logic_vector(31 downto 0);
    signal CONCAT_u1_u11_1370_1370_delayed_7_0_1308 : std_logic_vector(10 downto 0);
    signal CONCAT_u24_u64_1364_1364_delayed_7_0_1300 : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u106_1273_wire : std_logic_vector(105 downto 0);
    signal CONCAT_u32_u42_1018_wire : std_logic_vector(41 downto 0);
    signal CONCAT_u32_u64_1270_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1313_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u64_u74_1272_wire : std_logic_vector(73 downto 0);
    signal CONCAT_u64_u75_1315_wire : std_logic_vector(74 downto 0);
    signal CONCAT_u8_u16_1255_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_1258_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_1293_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u40_1298_wire : std_logic_vector(39 downto 0);
    signal EQ_u8_u1_1321_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1329_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1333_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1350_1350_delayed_7_0_1280 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1376_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_929_wire : std_logic_vector(0 downto 0);
    signal MUX_1019_wire : std_logic_vector(41 downto 0);
    signal MUX_1028_wire : std_logic_vector(41 downto 0);
    signal MUX_1117_wire : std_logic_vector(31 downto 0);
    signal MUX_1126_wire : std_logic_vector(31 downto 0);
    signal MUX_1336_wire : std_logic_vector(31 downto 0);
    signal MUX_1351_wire : std_logic_vector(31 downto 0);
    signal MUX_1352_wire : std_logic_vector(31 downto 0);
    signal MUX_996_wire : std_logic_vector(9 downto 0);
    signal NOT_u1_u1_1377_wire : std_logic_vector(0 downto 0);
    signal R_HALT_1375_wire_constant : std_logic_vector(7 downto 0);
    signal R_LOAD_1278_wire_constant : std_logic_vector(7 downto 0);
    signal R_one_10_935_wire_constant : std_logic_vector(9 downto 0);
    signal R_one_8_928_wire_constant : std_logic_vector(7 downto 0);
    signal R_read_signal_985_wire_constant : std_logic_vector(0 downto 0);
    signal R_zero_106_1266_wire_constant : std_logic_vector(105 downto 0);
    signal R_zero_10_992_wire_constant : std_logic_vector(9 downto 0);
    signal R_zero_139_1139_wire_constant : std_logic_vector(138 downto 0);
    signal R_zero_32_987_wire_constant : std_logic_vector(31 downto 0);
    signal R_zero_42_1013_wire_constant : std_logic_vector(41 downto 0);
    signal R_zero_42_1024_wire_constant : std_logic_vector(41 downto 0);
    signal cmd_925 : std_logic_vector(7 downto 0);
    signal dcache_actions_984 : std_logic_vector(2 downto 0);
    signal dcache_data_to_be_written_to_reg_1289 : std_logic_vector(31 downto 0);
    signal dcache_exec_result_1074 : std_logic_vector(31 downto 0);
    signal dcache_exec_result_1352_delayed_7_0_1283 : std_logic_vector(31 downto 0);
    signal dcache_isBranch_1078 : std_logic_vector(0 downto 0);
    signal dcache_opcode_1050 : std_logic_vector(7 downto 0);
    signal dcache_pc_1082 : std_logic_vector(9 downto 0);
    signal dcache_rd1_1066 : std_logic_vector(31 downto 0);
    signal dcache_rd2_1070 : std_logic_vector(31 downto 0);
    signal dcache_rd2_1365_delayed_7_0_1303 : std_logic_vector(31 downto 0);
    signal dcache_rd_1062 : std_logic_vector(7 downto 0);
    signal dcache_rs1_imm_1054 : std_logic_vector(7 downto 0);
    signal dcache_rs2_1058 : std_logic_vector(7 downto 0);
    signal dcache_state_953 : std_logic_vector(138 downto 0);
    signal dcache_to_ex_addr_32_1338 : std_logic_vector(31 downto 0);
    signal dcache_to_ex_rs1_imm_1098 : std_logic_vector(0 downto 0);
    signal dcache_to_ex_rs2_1102 : std_logic_vector(0 downto 0);
    signal ex_Unconditional_JUMP_984 : std_logic_vector(0 downto 0);
    signal final_memAddr_32_1166 : std_logic_vector(31 downto 0);
    signal final_rd1_1236 : std_logic_vector(31 downto 0);
    signal final_rd2_1248 : std_logic_vector(31 downto 0);
    signal flush_dcache_1221_delayed_4_0_1136 : std_logic_vector(0 downto 0);
    signal flush_dcache_984 : std_logic_vector(0 downto 0);
    signal flush_icache_984 : std_logic_vector(0 downto 0);
    signal flush_idecode_1058_delayed_7_0_1001 : std_logic_vector(0 downto 0);
    signal flush_idecode_984 : std_logic_vector(0 downto 0);
    signal flush_iexec_1330_delayed_7_0_1251 : std_logic_vector(0 downto 0);
    signal flush_iexec_984 : std_logic_vector(0 downto 0);
    signal flush_ifetch_984 : std_logic_vector(0 downto 0);
    signal flush_reg_984 : std_logic_vector(0 downto 0);
    signal icache_actions_984 : std_logic_vector(9 downto 0);
    signal icache_instruction_989 : std_logic_vector(31 downto 0);
    signal icache_state_1063_delayed_7_0_1010 : std_logic_vector(9 downto 0);
    signal icache_state_937 : std_logic_vector(9 downto 0);
    signal idecode_actions_984 : std_logic_vector(41 downto 0);
    signal idecode_state_1061_delayed_7_0_1007 : std_logic_vector(41 downto 0);
    signal idecode_state_941 : std_logic_vector(41 downto 0);
    signal iexec_actions_984 : std_logic_vector(3 downto 0);
    signal iexec_rd1_1042 : std_logic_vector(31 downto 0);
    signal iexec_rd1_final_1119 : std_logic_vector(31 downto 0);
    signal iexec_rd2_1046 : std_logic_vector(31 downto 0);
    signal iexec_rd2_final_1128 : std_logic_vector(31 downto 0);
    signal iexec_rs1_imm_1038 : std_logic_vector(7 downto 0);
    signal iexec_state_949 : std_logic_vector(105 downto 0);
    signal ifetch_actions_984 : std_logic_vector(9 downto 0);
    signal ifetch_state_933 : std_logic_vector(9 downto 0);
    signal iregfile_actions_984 : std_logic_vector(4 downto 0);
    signal iregfile_pc_1034 : std_logic_vector(9 downto 0);
    signal iregfile_pc_1342_delayed_7_0_1263 : std_logic_vector(9 downto 0);
    signal iregfile_state_945 : std_logic_vector(41 downto 0);
    signal iretire_exec_result_memData_1094 : std_logic_vector(31 downto 0);
    signal iretire_opcode_1086 : std_logic_vector(7 downto 0);
    signal iretire_rd_1090 : std_logic_vector(7 downto 0);
    signal iretire_state_957 : std_logic_vector(138 downto 0);
    signal iretire_state_to_dcache_addr_1150 : std_logic_vector(0 downto 0);
    signal iretire_state_to_dcache_memData_1154 : std_logic_vector(0 downto 0);
    signal iretire_state_to_ex_rs1_imm_1106 : std_logic_vector(0 downto 0);
    signal iretire_state_to_ex_rs2_1110 : std_logic_vector(0 downto 0);
    signal iretire_state_to_rs1_imm_1191 : std_logic_vector(0 downto 0);
    signal iretire_state_to_rs1_imm_1318_delayed_7_0_1227 : std_logic_vector(0 downto 0);
    signal iretire_state_to_rs2_1195 : std_logic_vector(0 downto 0);
    signal iretire_state_to_rs2_1324_delayed_7_0_1239 : std_logic_vector(0 downto 0);
    signal iretire_to_dcache_addr_32_1325 : std_logic_vector(31 downto 0);
    signal is_Branch_Hazard_984 : std_logic_vector(0 downto 0);
    signal konst_1348_wire_constant : std_logic_vector(9 downto 0);
    signal konst_939_wire_constant : std_logic_vector(9 downto 0);
    signal konst_943_wire_constant : std_logic_vector(41 downto 0);
    signal konst_947_wire_constant : std_logic_vector(41 downto 0);
    signal konst_951_wire_constant : std_logic_vector(105 downto 0);
    signal konst_955_wire_constant : std_logic_vector(138 downto 0);
    signal konst_959_wire_constant : std_logic_vector(138 downto 0);
    signal memAddr_1170 : std_logic_vector(9 downto 0);
    signal memReadData_1175 : std_logic_vector(31 downto 0);
    signal memWriteData_1160 : std_logic_vector(31 downto 0);
    signal memWrite_1146 : std_logic_vector(0 downto 0);
    signal n_dcache_state_1142 : std_logic_vector(138 downto 0);
    signal n_dcache_state_1142_956_buffered : std_logic_vector(138 downto 0);
    signal n_dcache_state_from_exec_1133 : std_logic_vector(138 downto 0);
    signal n_iRetire_state_1317 : std_logic_vector(138 downto 0);
    signal n_iRetire_state_1317_960_buffered : std_logic_vector(138 downto 0);
    signal n_icache_state_998 : std_logic_vector(9 downto 0);
    signal n_icache_state_998_940_buffered : std_logic_vector(9 downto 0);
    signal n_idecode_state_1021 : std_logic_vector(41 downto 0);
    signal n_idecode_state_1021_944_buffered : std_logic_vector(41 downto 0);
    signal n_iexec_state_1275 : std_logic_vector(105 downto 0);
    signal n_iexec_state_1275_952_buffered : std_logic_vector(105 downto 0);
    signal n_iregfile_state_1030 : std_logic_vector(41 downto 0);
    signal n_iregfile_state_1030_948_buffered : std_logic_vector(41 downto 0);
    signal next_ifetch_state_1358 : std_logic_vector(9 downto 0);
    signal next_ifetch_state_1358_936_buffered : std_logic_vector(9 downto 0);
    signal next_ifetch_state_32_1354 : std_logic_vector(31 downto 0);
    signal reg_d1_1224 : std_logic_vector(31 downto 0);
    signal reg_d2_1224 : std_logic_vector(31 downto 0);
    signal reg_data_to_be_written_1214 : std_logic_vector(31 downto 0);
    signal reg_data_to_be_written_1319_delayed_7_0_1230 : std_logic_vector(31 downto 0);
    signal reg_data_to_be_written_1325_delayed_7_0_1242 : std_logic_vector(31 downto 0);
    signal reg_opcode_1199 : std_logic_vector(7 downto 0);
    signal reg_rd_1211 : std_logic_vector(7 downto 0);
    signal reg_rs1_imm_1203 : std_logic_vector(7 downto 0);
    signal reg_rs2_1207 : std_logic_vector(7 downto 0);
    signal reg_valid_read1_1179 : std_logic_vector(0 downto 0);
    signal reg_valid_read2_1183 : std_logic_vector(0 downto 0);
    signal reg_valid_write_1187 : std_logic_vector(0 downto 0);
    signal stall_first_4_1060_delayed_7_0_1004 : std_logic_vector(0 downto 0);
    signal stall_first_4_984 : std_logic_vector(0 downto 0);
    signal type_cast_1346_wire : std_logic_vector(31 downto 0);
    signal type_cast_1350_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_HALT_1375_wire_constant <= "00000001";
    R_LOAD_1278_wire_constant <= "00000011";
    R_one_10_935_wire_constant <= "0000000001";
    R_one_8_928_wire_constant <= "00000001";
    R_read_signal_985_wire_constant <= "1";
    R_zero_106_1266_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    R_zero_10_992_wire_constant <= "0000000000";
    R_zero_139_1139_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    R_zero_32_987_wire_constant <= "00000000000000000000000000000000";
    R_zero_42_1013_wire_constant <= "000000000000000000000000000000000000000000";
    R_zero_42_1024_wire_constant <= "000000000000000000000000000000000000000000";
    konst_1348_wire_constant <= "0000000001";
    konst_939_wire_constant <= "0000000000";
    konst_943_wire_constant <= "000000000000000000000000000000000000000000";
    konst_947_wire_constant <= "000000000000000000000000000000000000000000";
    konst_951_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    konst_955_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    konst_959_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    -- logger for phi phi_stmt_933
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_933_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_933:input-0 R_one_10_935_wire_constant= " & Convert_SLV_To_Hex_String(R_one_10_935_wire_constant));
          --
        end if;
        if phi_stmt_933_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_933:input-1 next_ifetch_state_1358_936_buffered= " & Convert_SLV_To_Hex_String(next_ifetch_state_1358_936_buffered));
          --
        end if;
        if phi_stmt_933_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:processor_daemon:DP:phi_stmt_933:sample-completed");
          --
        end if;
        if phi_stmt_933_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:processor_daemon:DP:phi_stmt_933:output ifetch_state_933= " & Convert_SLV_To_Hex_String(ifetch_state_933));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_933: Block -- phi operator 
      signal idata: std_logic_vector(19 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_one_10_935_wire_constant & next_ifetch_state_1358_936_buffered;
      req <= phi_stmt_933_req_0 & phi_stmt_933_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_933",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 10) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_933_ack_0,
          idata => idata,
          odata => ifetch_state_933,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_933
    -- logger for phi phi_stmt_937
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_937_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_937:input-0 konst_939_wire_constant= " & Convert_SLV_To_Hex_String(konst_939_wire_constant));
          --
        end if;
        if phi_stmt_937_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_937:input-1 n_icache_state_998_940_buffered= " & Convert_SLV_To_Hex_String(n_icache_state_998_940_buffered));
          --
        end if;
        if phi_stmt_937_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:processor_daemon:DP:phi_stmt_937:sample-completed");
          --
        end if;
        if phi_stmt_937_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:processor_daemon:DP:phi_stmt_937:output icache_state_937= " & Convert_SLV_To_Hex_String(icache_state_937));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_937: Block -- phi operator 
      signal idata: std_logic_vector(19 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_939_wire_constant & n_icache_state_998_940_buffered;
      req <= phi_stmt_937_req_0 & phi_stmt_937_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_937",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 10) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_937_ack_0,
          idata => idata,
          odata => icache_state_937,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_937
    -- logger for phi phi_stmt_941
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_941_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_941:input-0 konst_943_wire_constant= " & Convert_SLV_To_Hex_String(konst_943_wire_constant));
          --
        end if;
        if phi_stmt_941_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_941:input-1 n_idecode_state_1021_944_buffered= " & Convert_SLV_To_Hex_String(n_idecode_state_1021_944_buffered));
          --
        end if;
        if phi_stmt_941_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:processor_daemon:DP:phi_stmt_941:sample-completed");
          --
        end if;
        if phi_stmt_941_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:processor_daemon:DP:phi_stmt_941:output idecode_state_941= " & Convert_SLV_To_Hex_String(idecode_state_941));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_941: Block -- phi operator 
      signal idata: std_logic_vector(83 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_943_wire_constant & n_idecode_state_1021_944_buffered;
      req <= phi_stmt_941_req_0 & phi_stmt_941_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_941",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 42) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_941_ack_0,
          idata => idata,
          odata => idecode_state_941,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_941
    -- logger for phi phi_stmt_945
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_945_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_945:input-0 konst_947_wire_constant= " & Convert_SLV_To_Hex_String(konst_947_wire_constant));
          --
        end if;
        if phi_stmt_945_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_945:input-1 n_iregfile_state_1030_948_buffered= " & Convert_SLV_To_Hex_String(n_iregfile_state_1030_948_buffered));
          --
        end if;
        if phi_stmt_945_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:processor_daemon:DP:phi_stmt_945:sample-completed");
          --
        end if;
        if phi_stmt_945_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:processor_daemon:DP:phi_stmt_945:output iregfile_state_945= " & Convert_SLV_To_Hex_String(iregfile_state_945));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_945: Block -- phi operator 
      signal idata: std_logic_vector(83 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_947_wire_constant & n_iregfile_state_1030_948_buffered;
      req <= phi_stmt_945_req_0 & phi_stmt_945_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_945",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 42) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_945_ack_0,
          idata => idata,
          odata => iregfile_state_945,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_945
    -- logger for phi phi_stmt_949
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_949_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_949:input-0 konst_951_wire_constant= " & Convert_SLV_To_Hex_String(konst_951_wire_constant));
          --
        end if;
        if phi_stmt_949_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_949:input-1 n_iexec_state_1275_952_buffered= " & Convert_SLV_To_Hex_String(n_iexec_state_1275_952_buffered));
          --
        end if;
        if phi_stmt_949_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:processor_daemon:DP:phi_stmt_949:sample-completed");
          --
        end if;
        if phi_stmt_949_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:processor_daemon:DP:phi_stmt_949:output iexec_state_949= " & Convert_SLV_To_Hex_String(iexec_state_949));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_949: Block -- phi operator 
      signal idata: std_logic_vector(211 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_951_wire_constant & n_iexec_state_1275_952_buffered;
      req <= phi_stmt_949_req_0 & phi_stmt_949_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_949",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 106) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_949_ack_0,
          idata => idata,
          odata => iexec_state_949,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_949
    -- logger for phi phi_stmt_953
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_953_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_953:input-0 konst_955_wire_constant= " & Convert_SLV_To_Hex_String(konst_955_wire_constant));
          --
        end if;
        if phi_stmt_953_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_953:input-1 n_dcache_state_1142_956_buffered= " & Convert_SLV_To_Hex_String(n_dcache_state_1142_956_buffered));
          --
        end if;
        if phi_stmt_953_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:processor_daemon:DP:phi_stmt_953:sample-completed");
          --
        end if;
        if phi_stmt_953_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:processor_daemon:DP:phi_stmt_953:output dcache_state_953= " & Convert_SLV_To_Hex_String(dcache_state_953));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_953: Block -- phi operator 
      signal idata: std_logic_vector(277 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_955_wire_constant & n_dcache_state_1142_956_buffered;
      req <= phi_stmt_953_req_0 & phi_stmt_953_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_953",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 139) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_953_ack_0,
          idata => idata,
          odata => dcache_state_953,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_953
    -- logger for phi phi_stmt_957
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_957_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_957:input-0 konst_959_wire_constant= " & Convert_SLV_To_Hex_String(konst_959_wire_constant));
          --
        end if;
        if phi_stmt_957_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:processor_daemon:DP:phi_stmt_957:input-1 n_iRetire_state_1317_960_buffered= " & Convert_SLV_To_Hex_String(n_iRetire_state_1317_960_buffered));
          --
        end if;
        if phi_stmt_957_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:processor_daemon:DP:phi_stmt_957:sample-completed");
          --
        end if;
        if phi_stmt_957_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:processor_daemon:DP:phi_stmt_957:output iretire_state_957= " & Convert_SLV_To_Hex_String(iretire_state_957));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_957: Block -- phi operator 
      signal idata: std_logic_vector(277 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_959_wire_constant & n_iRetire_state_1317_960_buffered;
      req <= phi_stmt_957_req_0 & phi_stmt_957_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_957",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 139) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_957_ack_0,
          idata => idata,
          odata => iretire_state_957,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_957
    -- logger for split-operator MUX_1019_inst flow-through 
    process(MUX_1019_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1019_inst:flowthrough inputs: " & " stall_first_4_1060_delayed_7_0_1004 = "& Convert_SLV_To_Hex_String(stall_first_4_1060_delayed_7_0_1004) & " idecode_state_1061_delayed_7_0_1007 = "& Convert_SLV_To_Hex_String(idecode_state_1061_delayed_7_0_1007) & " CONCAT_u32_u42_1018_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u42_1018_wire) & " outputs:" & " MUX_1019_wire= "  & Convert_SLV_To_Hex_String(MUX_1019_wire));
      --
    end process; 
    -- flow-through select operator MUX_1019_inst
    MUX_1019_wire <= idecode_state_1061_delayed_7_0_1007 when (stall_first_4_1060_delayed_7_0_1004(0) /=  '0') else CONCAT_u32_u42_1018_wire;
    -- logger for split-operator MUX_1020_inst flow-through 
    process(n_idecode_state_1021) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1020_inst:flowthrough inputs: " & " flush_idecode_1058_delayed_7_0_1001 = "& Convert_SLV_To_Hex_String(flush_idecode_1058_delayed_7_0_1001) & " R_zero_42_1013_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_42_1013_wire_constant) & " MUX_1019_wire = "& Convert_SLV_To_Hex_String(MUX_1019_wire) & " outputs:" & " n_idecode_state_1021= "  & Convert_SLV_To_Hex_String(n_idecode_state_1021));
      --
    end process; 
    -- flow-through select operator MUX_1020_inst
    n_idecode_state_1021 <= R_zero_42_1013_wire_constant when (flush_idecode_1058_delayed_7_0_1001(0) /=  '0') else MUX_1019_wire;
    -- logger for split-operator MUX_1028_inst flow-through 
    process(MUX_1028_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1028_inst:flowthrough inputs: " & " stall_first_4_984 = "& Convert_SLV_To_Hex_String(stall_first_4_984) & " iregfile_state_945 = "& Convert_SLV_To_Hex_String(iregfile_state_945) & " idecode_state_941 = "& Convert_SLV_To_Hex_String(idecode_state_941) & " outputs:" & " MUX_1028_wire= "  & Convert_SLV_To_Hex_String(MUX_1028_wire));
      --
    end process; 
    -- flow-through select operator MUX_1028_inst
    MUX_1028_wire <= iregfile_state_945 when (stall_first_4_984(0) /=  '0') else idecode_state_941;
    -- logger for split-operator MUX_1029_inst flow-through 
    process(n_iregfile_state_1030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1029_inst:flowthrough inputs: " & " flush_reg_984 = "& Convert_SLV_To_Hex_String(flush_reg_984) & " R_zero_42_1024_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_42_1024_wire_constant) & " MUX_1028_wire = "& Convert_SLV_To_Hex_String(MUX_1028_wire) & " outputs:" & " n_iregfile_state_1030= "  & Convert_SLV_To_Hex_String(n_iregfile_state_1030));
      --
    end process; 
    -- flow-through select operator MUX_1029_inst
    n_iregfile_state_1030 <= R_zero_42_1024_wire_constant when (flush_reg_984(0) /=  '0') else MUX_1028_wire;
    -- logger for split-operator MUX_1117_inst flow-through 
    process(MUX_1117_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1117_inst:flowthrough inputs: " & " iretire_state_to_ex_rs1_imm_1106 = "& Convert_SLV_To_Hex_String(iretire_state_to_ex_rs1_imm_1106) & " iretire_exec_result_memData_1094 = "& Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094) & " iexec_rd1_1042 = "& Convert_SLV_To_Hex_String(iexec_rd1_1042) & " outputs:" & " MUX_1117_wire= "  & Convert_SLV_To_Hex_String(MUX_1117_wire));
      --
    end process; 
    -- flow-through select operator MUX_1117_inst
    MUX_1117_wire <= iretire_exec_result_memData_1094 when (iretire_state_to_ex_rs1_imm_1106(0) /=  '0') else iexec_rd1_1042;
    -- logger for split-operator MUX_1118_inst flow-through 
    process(iexec_rd1_final_1119) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1118_inst:flowthrough inputs: " & " dcache_to_ex_rs1_imm_1098 = "& Convert_SLV_To_Hex_String(dcache_to_ex_rs1_imm_1098) & " dcache_exec_result_1074 = "& Convert_SLV_To_Hex_String(dcache_exec_result_1074) & " MUX_1117_wire = "& Convert_SLV_To_Hex_String(MUX_1117_wire) & " outputs:" & " iexec_rd1_final_1119= "  & Convert_SLV_To_Hex_String(iexec_rd1_final_1119));
      --
    end process; 
    -- flow-through select operator MUX_1118_inst
    iexec_rd1_final_1119 <= dcache_exec_result_1074 when (dcache_to_ex_rs1_imm_1098(0) /=  '0') else MUX_1117_wire;
    -- logger for split-operator MUX_1126_inst flow-through 
    process(MUX_1126_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1126_inst:flowthrough inputs: " & " iretire_state_to_ex_rs2_1110 = "& Convert_SLV_To_Hex_String(iretire_state_to_ex_rs2_1110) & " iretire_exec_result_memData_1094 = "& Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094) & " iexec_rd2_1046 = "& Convert_SLV_To_Hex_String(iexec_rd2_1046) & " outputs:" & " MUX_1126_wire= "  & Convert_SLV_To_Hex_String(MUX_1126_wire));
      --
    end process; 
    -- flow-through select operator MUX_1126_inst
    MUX_1126_wire <= iretire_exec_result_memData_1094 when (iretire_state_to_ex_rs2_1110(0) /=  '0') else iexec_rd2_1046;
    -- logger for split-operator MUX_1127_inst flow-through 
    process(iexec_rd2_final_1128) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1127_inst:flowthrough inputs: " & " dcache_to_ex_rs2_1102 = "& Convert_SLV_To_Hex_String(dcache_to_ex_rs2_1102) & " dcache_exec_result_1074 = "& Convert_SLV_To_Hex_String(dcache_exec_result_1074) & " MUX_1126_wire = "& Convert_SLV_To_Hex_String(MUX_1126_wire) & " outputs:" & " iexec_rd2_final_1128= "  & Convert_SLV_To_Hex_String(iexec_rd2_final_1128));
      --
    end process; 
    -- flow-through select operator MUX_1127_inst
    iexec_rd2_final_1128 <= dcache_exec_result_1074 when (dcache_to_ex_rs2_1102(0) /=  '0') else MUX_1126_wire;
    -- logger for split-operator MUX_1141_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_1141_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1141_inst:started:   inputs: " & " flush_dcache_1221_delayed_4_0_1136 = "& Convert_SLV_To_Hex_String(flush_dcache_1221_delayed_4_0_1136) & " R_zero_139_1139_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_139_1139_wire_constant) & " n_dcache_state_from_exec_1133 = "& Convert_SLV_To_Hex_String(n_dcache_state_from_exec_1133));
          --
        end if; 
        if MUX_1141_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1141_inst:finished:  outputs: " & " n_dcache_state_1142= "  & Convert_SLV_To_Hex_String(n_dcache_state_1142));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_1141_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1141_inst_req_0;
      MUX_1141_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1141_inst_req_1;
      MUX_1141_inst_ack_1<= update_ack(0);
      MUX_1141_inst: SelectSplitProtocol generic map(name => "MUX_1141_inst", data_width => 139, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => R_zero_139_1139_wire_constant, y => n_dcache_state_from_exec_1133, sel => flush_dcache_1221_delayed_4_0_1136, z => n_dcache_state_1142, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator MUX_1159_inst flow-through 
    process(memWriteData_1160) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1159_inst:flowthrough inputs: " & " iretire_state_to_dcache_memData_1154 = "& Convert_SLV_To_Hex_String(iretire_state_to_dcache_memData_1154) & " iretire_exec_result_memData_1094 = "& Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094) & " dcache_rd2_1070 = "& Convert_SLV_To_Hex_String(dcache_rd2_1070) & " outputs:" & " memWriteData_1160= "  & Convert_SLV_To_Hex_String(memWriteData_1160));
      --
    end process; 
    -- flow-through select operator MUX_1159_inst
    memWriteData_1160 <= iretire_exec_result_memData_1094 when (iretire_state_to_dcache_memData_1154(0) /=  '0') else dcache_rd2_1070;
    -- logger for split-operator MUX_1165_inst flow-through 
    process(final_memAddr_32_1166) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1165_inst:flowthrough inputs: " & " iretire_state_to_dcache_addr_1150 = "& Convert_SLV_To_Hex_String(iretire_state_to_dcache_addr_1150) & " iretire_exec_result_memData_1094 = "& Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094) & " dcache_rd1_1066 = "& Convert_SLV_To_Hex_String(dcache_rd1_1066) & " outputs:" & " final_memAddr_32_1166= "  & Convert_SLV_To_Hex_String(final_memAddr_32_1166));
      --
    end process; 
    -- flow-through select operator MUX_1165_inst
    final_memAddr_32_1166 <= iretire_exec_result_memData_1094 when (iretire_state_to_dcache_addr_1150(0) /=  '0') else dcache_rd1_1066;
    -- logger for split-operator MUX_1235_inst flow-through 
    process(final_rd1_1236) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1235_inst:flowthrough inputs: " & " iretire_state_to_rs1_imm_1318_delayed_7_0_1227 = "& Convert_SLV_To_Hex_String(iretire_state_to_rs1_imm_1318_delayed_7_0_1227) & " reg_data_to_be_written_1319_delayed_7_0_1230 = "& Convert_SLV_To_Hex_String(reg_data_to_be_written_1319_delayed_7_0_1230) & " reg_d1_1224 = "& Convert_SLV_To_Hex_String(reg_d1_1224) & " outputs:" & " final_rd1_1236= "  & Convert_SLV_To_Hex_String(final_rd1_1236));
      --
    end process; 
    -- flow-through select operator MUX_1235_inst
    final_rd1_1236 <= reg_data_to_be_written_1319_delayed_7_0_1230 when (iretire_state_to_rs1_imm_1318_delayed_7_0_1227(0) /=  '0') else reg_d1_1224;
    -- logger for split-operator MUX_1247_inst flow-through 
    process(final_rd2_1248) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1247_inst:flowthrough inputs: " & " iretire_state_to_rs2_1324_delayed_7_0_1239 = "& Convert_SLV_To_Hex_String(iretire_state_to_rs2_1324_delayed_7_0_1239) & " reg_data_to_be_written_1325_delayed_7_0_1242 = "& Convert_SLV_To_Hex_String(reg_data_to_be_written_1325_delayed_7_0_1242) & " reg_d2_1224 = "& Convert_SLV_To_Hex_String(reg_d2_1224) & " outputs:" & " final_rd2_1248= "  & Convert_SLV_To_Hex_String(final_rd2_1248));
      --
    end process; 
    -- flow-through select operator MUX_1247_inst
    final_rd2_1248 <= reg_data_to_be_written_1325_delayed_7_0_1242 when (iretire_state_to_rs2_1324_delayed_7_0_1239(0) /=  '0') else reg_d2_1224;
    -- logger for split-operator MUX_1274_inst flow-through 
    process(n_iexec_state_1275) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1274_inst:flowthrough inputs: " & " flush_iexec_1330_delayed_7_0_1251 = "& Convert_SLV_To_Hex_String(flush_iexec_1330_delayed_7_0_1251) & " R_zero_106_1266_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_106_1266_wire_constant) & " CONCAT_u32_u106_1273_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u106_1273_wire) & " outputs:" & " n_iexec_state_1275= "  & Convert_SLV_To_Hex_String(n_iexec_state_1275));
      --
    end process; 
    -- flow-through select operator MUX_1274_inst
    n_iexec_state_1275 <= R_zero_106_1266_wire_constant when (flush_iexec_1330_delayed_7_0_1251(0) /=  '0') else CONCAT_u32_u106_1273_wire;
    -- logger for split-operator MUX_1288_inst flow-through 
    process(dcache_data_to_be_written_to_reg_1289) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1288_inst:flowthrough inputs: " & " EQ_u8_u1_1350_1350_delayed_7_0_1280 = "& Convert_SLV_To_Hex_String(EQ_u8_u1_1350_1350_delayed_7_0_1280) & " memReadData_1175 = "& Convert_SLV_To_Hex_String(memReadData_1175) & " dcache_exec_result_1352_delayed_7_0_1283 = "& Convert_SLV_To_Hex_String(dcache_exec_result_1352_delayed_7_0_1283) & " outputs:" & " dcache_data_to_be_written_to_reg_1289= "  & Convert_SLV_To_Hex_String(dcache_data_to_be_written_to_reg_1289));
      --
    end process; 
    -- flow-through select operator MUX_1288_inst
    dcache_data_to_be_written_to_reg_1289 <= memReadData_1175 when (EQ_u8_u1_1350_1350_delayed_7_0_1280(0) /=  '0') else dcache_exec_result_1352_delayed_7_0_1283;
    -- logger for split-operator MUX_1324_inst flow-through 
    process(iretire_to_dcache_addr_32_1325) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1324_inst:flowthrough inputs: " & " EQ_u8_u1_1321_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_1321_wire) & " iretire_exec_result_memData_1094 = "& Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094) & " dcache_rd2_1070 = "& Convert_SLV_To_Hex_String(dcache_rd2_1070) & " outputs:" & " iretire_to_dcache_addr_32_1325= "  & Convert_SLV_To_Hex_String(iretire_to_dcache_addr_32_1325));
      --
    end process; 
    -- flow-through select operator MUX_1324_inst
    iretire_to_dcache_addr_32_1325 <= iretire_exec_result_memData_1094 when (EQ_u8_u1_1321_wire(0) /=  '0') else dcache_rd2_1070;
    -- logger for split-operator MUX_1336_inst flow-through 
    process(MUX_1336_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1336_inst:flowthrough inputs: " & " EQ_u8_u1_1333_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_1333_wire) & " iretire_exec_result_memData_1094 = "& Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094) & " iexec_rd1_1042 = "& Convert_SLV_To_Hex_String(iexec_rd1_1042) & " outputs:" & " MUX_1336_wire= "  & Convert_SLV_To_Hex_String(MUX_1336_wire));
      --
    end process; 
    -- flow-through select operator MUX_1336_inst
    MUX_1336_wire <= iretire_exec_result_memData_1094 when (EQ_u8_u1_1333_wire(0) /=  '0') else iexec_rd1_1042;
    -- logger for split-operator MUX_1337_inst flow-through 
    process(dcache_to_ex_addr_32_1338) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1337_inst:flowthrough inputs: " & " EQ_u8_u1_1329_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_1329_wire) & " dcache_exec_result_1074 = "& Convert_SLV_To_Hex_String(dcache_exec_result_1074) & " MUX_1336_wire = "& Convert_SLV_To_Hex_String(MUX_1336_wire) & " outputs:" & " dcache_to_ex_addr_32_1338= "  & Convert_SLV_To_Hex_String(dcache_to_ex_addr_32_1338));
      --
    end process; 
    -- flow-through select operator MUX_1337_inst
    dcache_to_ex_addr_32_1338 <= dcache_exec_result_1074 when (EQ_u8_u1_1329_wire(0) /=  '0') else MUX_1336_wire;
    -- logger for split-operator MUX_1351_inst flow-through 
    process(MUX_1351_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1351_inst:flowthrough inputs: " & " stall_first_4_984 = "& Convert_SLV_To_Hex_String(stall_first_4_984) & " type_cast_1346_wire = "& Convert_SLV_To_Hex_String(type_cast_1346_wire) & " type_cast_1350_wire = "& Convert_SLV_To_Hex_String(type_cast_1350_wire) & " outputs:" & " MUX_1351_wire= "  & Convert_SLV_To_Hex_String(MUX_1351_wire));
      --
    end process; 
    -- flow-through select operator MUX_1351_inst
    MUX_1351_wire <= type_cast_1346_wire when (stall_first_4_984(0) /=  '0') else type_cast_1350_wire;
    -- logger for split-operator MUX_1352_inst flow-through 
    process(MUX_1352_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1352_inst:flowthrough inputs: " & " ex_Unconditional_JUMP_984 = "& Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_984) & " dcache_to_ex_addr_32_1338 = "& Convert_SLV_To_Hex_String(dcache_to_ex_addr_32_1338) & " MUX_1351_wire = "& Convert_SLV_To_Hex_String(MUX_1351_wire) & " outputs:" & " MUX_1352_wire= "  & Convert_SLV_To_Hex_String(MUX_1352_wire));
      --
    end process; 
    -- flow-through select operator MUX_1352_inst
    MUX_1352_wire <= dcache_to_ex_addr_32_1338 when (ex_Unconditional_JUMP_984(0) /=  '0') else MUX_1351_wire;
    -- logger for split-operator MUX_1353_inst flow-through 
    process(next_ifetch_state_32_1354) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_1353_inst:flowthrough inputs: " & " is_Branch_Hazard_984 = "& Convert_SLV_To_Hex_String(is_Branch_Hazard_984) & " iretire_to_dcache_addr_32_1325 = "& Convert_SLV_To_Hex_String(iretire_to_dcache_addr_32_1325) & " MUX_1352_wire = "& Convert_SLV_To_Hex_String(MUX_1352_wire) & " outputs:" & " next_ifetch_state_32_1354= "  & Convert_SLV_To_Hex_String(next_ifetch_state_32_1354));
      --
    end process; 
    -- flow-through select operator MUX_1353_inst
    next_ifetch_state_32_1354 <= iretire_to_dcache_addr_32_1325 when (is_Branch_Hazard_984(0) /=  '0') else MUX_1352_wire;
    -- logger for split-operator MUX_996_inst flow-through 
    process(MUX_996_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_996_inst:flowthrough inputs: " & " stall_first_4_984 = "& Convert_SLV_To_Hex_String(stall_first_4_984) & " icache_state_937 = "& Convert_SLV_To_Hex_String(icache_state_937) & " ifetch_state_933 = "& Convert_SLV_To_Hex_String(ifetch_state_933) & " outputs:" & " MUX_996_wire= "  & Convert_SLV_To_Hex_String(MUX_996_wire));
      --
    end process; 
    -- flow-through select operator MUX_996_inst
    MUX_996_wire <= icache_state_937 when (stall_first_4_984(0) /=  '0') else ifetch_state_933;
    -- logger for split-operator MUX_997_inst flow-through 
    process(n_icache_state_998) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:MUX_997_inst:flowthrough inputs: " & " flush_icache_984 = "& Convert_SLV_To_Hex_String(flush_icache_984) & " R_zero_10_992_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_10_992_wire_constant) & " MUX_996_wire = "& Convert_SLV_To_Hex_String(MUX_996_wire) & " outputs:" & " n_icache_state_998= "  & Convert_SLV_To_Hex_String(n_icache_state_998));
      --
    end process; 
    -- flow-through select operator MUX_997_inst
    n_icache_state_998 <= R_zero_10_992_wire_constant when (flush_icache_984(0) /=  '0') else MUX_996_wire;
    -- logger for split-operator slice_1033_inst flow-through 
    process(iregfile_pc_1034) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1033_inst:flowthrough inputs: " & " iregfile_state_945 = "& Convert_SLV_To_Hex_String(iregfile_state_945) & " outputs:" & " iregfile_pc_1034= "  & Convert_SLV_To_Hex_String(iregfile_pc_1034));
      --
    end process; 
    -- flow-through slice operator slice_1033_inst
    iregfile_pc_1034 <= iregfile_state_945(9 downto 0);
    -- logger for split-operator slice_1037_inst flow-through 
    process(iexec_rs1_imm_1038) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1037_inst:flowthrough inputs: " & " iexec_state_949 = "& Convert_SLV_To_Hex_String(iexec_state_949) & " outputs:" & " iexec_rs1_imm_1038= "  & Convert_SLV_To_Hex_String(iexec_rs1_imm_1038));
      --
    end process; 
    -- flow-through slice operator slice_1037_inst
    iexec_rs1_imm_1038 <= iexec_state_949(97 downto 90);
    -- logger for split-operator slice_1041_inst flow-through 
    process(iexec_rd1_1042) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1041_inst:flowthrough inputs: " & " iexec_state_949 = "& Convert_SLV_To_Hex_String(iexec_state_949) & " outputs:" & " iexec_rd1_1042= "  & Convert_SLV_To_Hex_String(iexec_rd1_1042));
      --
    end process; 
    -- flow-through slice operator slice_1041_inst
    iexec_rd1_1042 <= iexec_state_949(73 downto 42);
    -- logger for split-operator slice_1045_inst flow-through 
    process(iexec_rd2_1046) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1045_inst:flowthrough inputs: " & " iexec_state_949 = "& Convert_SLV_To_Hex_String(iexec_state_949) & " outputs:" & " iexec_rd2_1046= "  & Convert_SLV_To_Hex_String(iexec_rd2_1046));
      --
    end process; 
    -- flow-through slice operator slice_1045_inst
    iexec_rd2_1046 <= iexec_state_949(41 downto 10);
    -- logger for split-operator slice_1049_inst flow-through 
    process(dcache_opcode_1050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1049_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_opcode_1050= "  & Convert_SLV_To_Hex_String(dcache_opcode_1050));
      --
    end process; 
    -- flow-through slice operator slice_1049_inst
    dcache_opcode_1050 <= dcache_state_953(138 downto 131);
    -- logger for split-operator slice_1053_inst flow-through 
    process(dcache_rs1_imm_1054) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1053_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_rs1_imm_1054= "  & Convert_SLV_To_Hex_String(dcache_rs1_imm_1054));
      --
    end process; 
    -- flow-through slice operator slice_1053_inst
    dcache_rs1_imm_1054 <= dcache_state_953(130 downto 123);
    -- logger for split-operator slice_1057_inst flow-through 
    process(dcache_rs2_1058) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1057_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_rs2_1058= "  & Convert_SLV_To_Hex_String(dcache_rs2_1058));
      --
    end process; 
    -- flow-through slice operator slice_1057_inst
    dcache_rs2_1058 <= dcache_state_953(122 downto 115);
    -- logger for split-operator slice_1061_inst flow-through 
    process(dcache_rd_1062) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1061_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_rd_1062= "  & Convert_SLV_To_Hex_String(dcache_rd_1062));
      --
    end process; 
    -- flow-through slice operator slice_1061_inst
    dcache_rd_1062 <= dcache_state_953(114 downto 107);
    -- logger for split-operator slice_1065_inst flow-through 
    process(dcache_rd1_1066) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1065_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_rd1_1066= "  & Convert_SLV_To_Hex_String(dcache_rd1_1066));
      --
    end process; 
    -- flow-through slice operator slice_1065_inst
    dcache_rd1_1066 <= dcache_state_953(106 downto 75);
    -- logger for split-operator slice_1069_inst flow-through 
    process(dcache_rd2_1070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1069_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_rd2_1070= "  & Convert_SLV_To_Hex_String(dcache_rd2_1070));
      --
    end process; 
    -- flow-through slice operator slice_1069_inst
    dcache_rd2_1070 <= dcache_state_953(74 downto 43);
    -- logger for split-operator slice_1073_inst flow-through 
    process(dcache_exec_result_1074) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1073_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_exec_result_1074= "  & Convert_SLV_To_Hex_String(dcache_exec_result_1074));
      --
    end process; 
    -- flow-through slice operator slice_1073_inst
    dcache_exec_result_1074 <= dcache_state_953(42 downto 11);
    -- logger for split-operator slice_1077_inst flow-through 
    process(dcache_isBranch_1078) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1077_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_isBranch_1078= "  & Convert_SLV_To_Hex_String(dcache_isBranch_1078));
      --
    end process; 
    -- flow-through slice operator slice_1077_inst
    dcache_isBranch_1078 <= dcache_state_953(10 downto 10);
    -- logger for split-operator slice_1081_inst flow-through 
    process(dcache_pc_1082) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1081_inst:flowthrough inputs: " & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " outputs:" & " dcache_pc_1082= "  & Convert_SLV_To_Hex_String(dcache_pc_1082));
      --
    end process; 
    -- flow-through slice operator slice_1081_inst
    dcache_pc_1082 <= dcache_state_953(9 downto 0);
    -- logger for split-operator slice_1085_inst flow-through 
    process(iretire_opcode_1086) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1085_inst:flowthrough inputs: " & " iretire_state_957 = "& Convert_SLV_To_Hex_String(iretire_state_957) & " outputs:" & " iretire_opcode_1086= "  & Convert_SLV_To_Hex_String(iretire_opcode_1086));
      --
    end process; 
    -- flow-through slice operator slice_1085_inst
    iretire_opcode_1086 <= iretire_state_957(138 downto 131);
    -- logger for split-operator slice_1089_inst flow-through 
    process(iretire_rd_1090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1089_inst:flowthrough inputs: " & " iretire_state_957 = "& Convert_SLV_To_Hex_String(iretire_state_957) & " outputs:" & " iretire_rd_1090= "  & Convert_SLV_To_Hex_String(iretire_rd_1090));
      --
    end process; 
    -- flow-through slice operator slice_1089_inst
    iretire_rd_1090 <= iretire_state_957(114 downto 107);
    -- logger for split-operator slice_1093_inst flow-through 
    process(iretire_exec_result_memData_1094) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1093_inst:flowthrough inputs: " & " iretire_state_957 = "& Convert_SLV_To_Hex_String(iretire_state_957) & " outputs:" & " iretire_exec_result_memData_1094= "  & Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094));
      --
    end process; 
    -- flow-through slice operator slice_1093_inst
    iretire_exec_result_memData_1094 <= iretire_state_957(42 downto 11);
    -- logger for split-operator slice_1097_inst flow-through 
    process(dcache_to_ex_rs1_imm_1098) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1097_inst:flowthrough inputs: " & " iexec_actions_984 = "& Convert_SLV_To_Hex_String(iexec_actions_984) & " outputs:" & " dcache_to_ex_rs1_imm_1098= "  & Convert_SLV_To_Hex_String(dcache_to_ex_rs1_imm_1098));
      --
    end process; 
    -- flow-through slice operator slice_1097_inst
    dcache_to_ex_rs1_imm_1098 <= iexec_actions_984(3 downto 3);
    -- logger for split-operator slice_1101_inst flow-through 
    process(dcache_to_ex_rs2_1102) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1101_inst:flowthrough inputs: " & " iexec_actions_984 = "& Convert_SLV_To_Hex_String(iexec_actions_984) & " outputs:" & " dcache_to_ex_rs2_1102= "  & Convert_SLV_To_Hex_String(dcache_to_ex_rs2_1102));
      --
    end process; 
    -- flow-through slice operator slice_1101_inst
    dcache_to_ex_rs2_1102 <= iexec_actions_984(2 downto 2);
    -- logger for split-operator slice_1105_inst flow-through 
    process(iretire_state_to_ex_rs1_imm_1106) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1105_inst:flowthrough inputs: " & " iexec_actions_984 = "& Convert_SLV_To_Hex_String(iexec_actions_984) & " outputs:" & " iretire_state_to_ex_rs1_imm_1106= "  & Convert_SLV_To_Hex_String(iretire_state_to_ex_rs1_imm_1106));
      --
    end process; 
    -- flow-through slice operator slice_1105_inst
    iretire_state_to_ex_rs1_imm_1106 <= iexec_actions_984(1 downto 1);
    -- logger for split-operator slice_1109_inst flow-through 
    process(iretire_state_to_ex_rs2_1110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1109_inst:flowthrough inputs: " & " iexec_actions_984 = "& Convert_SLV_To_Hex_String(iexec_actions_984) & " outputs:" & " iretire_state_to_ex_rs2_1110= "  & Convert_SLV_To_Hex_String(iretire_state_to_ex_rs2_1110));
      --
    end process; 
    -- flow-through slice operator slice_1109_inst
    iretire_state_to_ex_rs2_1110 <= iexec_actions_984(0 downto 0);
    -- logger for split-operator slice_1145_inst flow-through 
    process(memWrite_1146) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1145_inst:flowthrough inputs: " & " dcache_actions_984 = "& Convert_SLV_To_Hex_String(dcache_actions_984) & " outputs:" & " memWrite_1146= "  & Convert_SLV_To_Hex_String(memWrite_1146));
      --
    end process; 
    -- flow-through slice operator slice_1145_inst
    memWrite_1146 <= dcache_actions_984(2 downto 2);
    -- logger for split-operator slice_1149_inst flow-through 
    process(iretire_state_to_dcache_addr_1150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1149_inst:flowthrough inputs: " & " dcache_actions_984 = "& Convert_SLV_To_Hex_String(dcache_actions_984) & " outputs:" & " iretire_state_to_dcache_addr_1150= "  & Convert_SLV_To_Hex_String(iretire_state_to_dcache_addr_1150));
      --
    end process; 
    -- flow-through slice operator slice_1149_inst
    iretire_state_to_dcache_addr_1150 <= dcache_actions_984(1 downto 1);
    -- logger for split-operator slice_1153_inst flow-through 
    process(iretire_state_to_dcache_memData_1154) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1153_inst:flowthrough inputs: " & " dcache_actions_984 = "& Convert_SLV_To_Hex_String(dcache_actions_984) & " outputs:" & " iretire_state_to_dcache_memData_1154= "  & Convert_SLV_To_Hex_String(iretire_state_to_dcache_memData_1154));
      --
    end process; 
    -- flow-through slice operator slice_1153_inst
    iretire_state_to_dcache_memData_1154 <= dcache_actions_984(0 downto 0);
    -- logger for split-operator slice_1169_inst flow-through 
    process(memAddr_1170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1169_inst:flowthrough inputs: " & " final_memAddr_32_1166 = "& Convert_SLV_To_Hex_String(final_memAddr_32_1166) & " outputs:" & " memAddr_1170= "  & Convert_SLV_To_Hex_String(memAddr_1170));
      --
    end process; 
    -- flow-through slice operator slice_1169_inst
    memAddr_1170 <= final_memAddr_32_1166(9 downto 0);
    -- logger for split-operator slice_1178_inst flow-through 
    process(reg_valid_read1_1179) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1178_inst:flowthrough inputs: " & " iregfile_actions_984 = "& Convert_SLV_To_Hex_String(iregfile_actions_984) & " outputs:" & " reg_valid_read1_1179= "  & Convert_SLV_To_Hex_String(reg_valid_read1_1179));
      --
    end process; 
    -- flow-through slice operator slice_1178_inst
    reg_valid_read1_1179 <= iregfile_actions_984(4 downto 4);
    -- logger for split-operator slice_1182_inst flow-through 
    process(reg_valid_read2_1183) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1182_inst:flowthrough inputs: " & " iregfile_actions_984 = "& Convert_SLV_To_Hex_String(iregfile_actions_984) & " outputs:" & " reg_valid_read2_1183= "  & Convert_SLV_To_Hex_String(reg_valid_read2_1183));
      --
    end process; 
    -- flow-through slice operator slice_1182_inst
    reg_valid_read2_1183 <= iregfile_actions_984(3 downto 3);
    -- logger for split-operator slice_1186_inst flow-through 
    process(reg_valid_write_1187) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1186_inst:flowthrough inputs: " & " iregfile_actions_984 = "& Convert_SLV_To_Hex_String(iregfile_actions_984) & " outputs:" & " reg_valid_write_1187= "  & Convert_SLV_To_Hex_String(reg_valid_write_1187));
      --
    end process; 
    -- flow-through slice operator slice_1186_inst
    reg_valid_write_1187 <= iregfile_actions_984(2 downto 2);
    -- logger for split-operator slice_1190_inst flow-through 
    process(iretire_state_to_rs1_imm_1191) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1190_inst:flowthrough inputs: " & " iregfile_actions_984 = "& Convert_SLV_To_Hex_String(iregfile_actions_984) & " outputs:" & " iretire_state_to_rs1_imm_1191= "  & Convert_SLV_To_Hex_String(iretire_state_to_rs1_imm_1191));
      --
    end process; 
    -- flow-through slice operator slice_1190_inst
    iretire_state_to_rs1_imm_1191 <= iregfile_actions_984(1 downto 1);
    -- logger for split-operator slice_1194_inst flow-through 
    process(iretire_state_to_rs2_1195) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1194_inst:flowthrough inputs: " & " iregfile_actions_984 = "& Convert_SLV_To_Hex_String(iregfile_actions_984) & " outputs:" & " iretire_state_to_rs2_1195= "  & Convert_SLV_To_Hex_String(iretire_state_to_rs2_1195));
      --
    end process; 
    -- flow-through slice operator slice_1194_inst
    iretire_state_to_rs2_1195 <= iregfile_actions_984(0 downto 0);
    -- logger for split-operator slice_1198_inst flow-through 
    process(reg_opcode_1199) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1198_inst:flowthrough inputs: " & " iregfile_state_945 = "& Convert_SLV_To_Hex_String(iregfile_state_945) & " outputs:" & " reg_opcode_1199= "  & Convert_SLV_To_Hex_String(reg_opcode_1199));
      --
    end process; 
    -- flow-through slice operator slice_1198_inst
    reg_opcode_1199 <= iregfile_state_945(41 downto 34);
    -- logger for split-operator slice_1202_inst flow-through 
    process(reg_rs1_imm_1203) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1202_inst:flowthrough inputs: " & " iregfile_state_945 = "& Convert_SLV_To_Hex_String(iregfile_state_945) & " outputs:" & " reg_rs1_imm_1203= "  & Convert_SLV_To_Hex_String(reg_rs1_imm_1203));
      --
    end process; 
    -- flow-through slice operator slice_1202_inst
    reg_rs1_imm_1203 <= iregfile_state_945(33 downto 26);
    -- logger for split-operator slice_1206_inst flow-through 
    process(reg_rs2_1207) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1206_inst:flowthrough inputs: " & " iregfile_state_945 = "& Convert_SLV_To_Hex_String(iregfile_state_945) & " outputs:" & " reg_rs2_1207= "  & Convert_SLV_To_Hex_String(reg_rs2_1207));
      --
    end process; 
    -- flow-through slice operator slice_1206_inst
    reg_rs2_1207 <= iregfile_state_945(25 downto 18);
    -- logger for split-operator slice_1210_inst flow-through 
    process(reg_rd_1211) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1210_inst:flowthrough inputs: " & " iregfile_state_945 = "& Convert_SLV_To_Hex_String(iregfile_state_945) & " outputs:" & " reg_rd_1211= "  & Convert_SLV_To_Hex_String(reg_rd_1211));
      --
    end process; 
    -- flow-through slice operator slice_1210_inst
    reg_rd_1211 <= iregfile_state_945(17 downto 10);
    -- logger for split-operator slice_1357_inst flow-through 
    process(next_ifetch_state_1358) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:slice_1357_inst:flowthrough inputs: " & " next_ifetch_state_32_1354 = "& Convert_SLV_To_Hex_String(next_ifetch_state_32_1354) & " outputs:" & " next_ifetch_state_1358= "  & Convert_SLV_To_Hex_String(next_ifetch_state_1358));
      --
    end process; 
    -- flow-through slice operator slice_1357_inst
    next_ifetch_state_1358 <= next_ifetch_state_32_1354(9 downto 0);
    -- logger for split-operator W_dcache_exec_result_1352_delayed_7_0_1281_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_dcache_exec_result_1352_delayed_7_0_1281_inst:started:   inputs: " & " dcache_exec_result_1074 = "& Convert_SLV_To_Hex_String(dcache_exec_result_1074));
          --
        end if; 
        if W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_dcache_exec_result_1352_delayed_7_0_1281_inst:finished:  outputs: " & " dcache_exec_result_1352_delayed_7_0_1283= "  & Convert_SLV_To_Hex_String(dcache_exec_result_1352_delayed_7_0_1283));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_dcache_exec_result_1352_delayed_7_0_1281_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_0;
      W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_0<= wack(0);
      rreq(0) <= W_dcache_exec_result_1352_delayed_7_0_1281_inst_req_1;
      W_dcache_exec_result_1352_delayed_7_0_1281_inst_ack_1<= rack(0);
      W_dcache_exec_result_1352_delayed_7_0_1281_inst : InterlockBuffer generic map ( -- 
        name => "W_dcache_exec_result_1352_delayed_7_0_1281_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => dcache_exec_result_1074,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => dcache_exec_result_1352_delayed_7_0_1283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_dcache_rd2_1365_delayed_7_0_1301_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_dcache_rd2_1365_delayed_7_0_1301_inst:started:   inputs: " & " dcache_rd2_1070 = "& Convert_SLV_To_Hex_String(dcache_rd2_1070));
          --
        end if; 
        if W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_dcache_rd2_1365_delayed_7_0_1301_inst:finished:  outputs: " & " dcache_rd2_1365_delayed_7_0_1303= "  & Convert_SLV_To_Hex_String(dcache_rd2_1365_delayed_7_0_1303));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_dcache_rd2_1365_delayed_7_0_1301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_dcache_rd2_1365_delayed_7_0_1301_inst_req_0;
      W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_0<= wack(0);
      rreq(0) <= W_dcache_rd2_1365_delayed_7_0_1301_inst_req_1;
      W_dcache_rd2_1365_delayed_7_0_1301_inst_ack_1<= rack(0);
      W_dcache_rd2_1365_delayed_7_0_1301_inst : InterlockBuffer generic map ( -- 
        name => "W_dcache_rd2_1365_delayed_7_0_1301_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => dcache_rd2_1070,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => dcache_rd2_1365_delayed_7_0_1303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_flush_dcache_1221_delayed_4_0_1134_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_flush_dcache_1221_delayed_4_0_1134_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_flush_dcache_1221_delayed_4_0_1134_inst:started:   inputs: " & " flush_dcache_984 = "& Convert_SLV_To_Hex_String(flush_dcache_984));
          --
        end if; 
        if W_flush_dcache_1221_delayed_4_0_1134_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_flush_dcache_1221_delayed_4_0_1134_inst:finished:  outputs: " & " flush_dcache_1221_delayed_4_0_1136= "  & Convert_SLV_To_Hex_String(flush_dcache_1221_delayed_4_0_1136));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_flush_dcache_1221_delayed_4_0_1134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_flush_dcache_1221_delayed_4_0_1134_inst_req_0;
      W_flush_dcache_1221_delayed_4_0_1134_inst_ack_0<= wack(0);
      rreq(0) <= W_flush_dcache_1221_delayed_4_0_1134_inst_req_1;
      W_flush_dcache_1221_delayed_4_0_1134_inst_ack_1<= rack(0);
      W_flush_dcache_1221_delayed_4_0_1134_inst : InterlockBuffer generic map ( -- 
        name => "W_flush_dcache_1221_delayed_4_0_1134_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => flush_dcache_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => flush_dcache_1221_delayed_4_0_1136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_flush_idecode_1058_delayed_7_0_999_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_flush_idecode_1058_delayed_7_0_999_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_flush_idecode_1058_delayed_7_0_999_inst:started:   inputs: " & " flush_idecode_984 = "& Convert_SLV_To_Hex_String(flush_idecode_984));
          --
        end if; 
        if W_flush_idecode_1058_delayed_7_0_999_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_flush_idecode_1058_delayed_7_0_999_inst:finished:  outputs: " & " flush_idecode_1058_delayed_7_0_1001= "  & Convert_SLV_To_Hex_String(flush_idecode_1058_delayed_7_0_1001));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_flush_idecode_1058_delayed_7_0_999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_flush_idecode_1058_delayed_7_0_999_inst_req_0;
      W_flush_idecode_1058_delayed_7_0_999_inst_ack_0<= wack(0);
      rreq(0) <= W_flush_idecode_1058_delayed_7_0_999_inst_req_1;
      W_flush_idecode_1058_delayed_7_0_999_inst_ack_1<= rack(0);
      W_flush_idecode_1058_delayed_7_0_999_inst : InterlockBuffer generic map ( -- 
        name => "W_flush_idecode_1058_delayed_7_0_999_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => flush_idecode_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => flush_idecode_1058_delayed_7_0_1001,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_flush_iexec_1330_delayed_7_0_1249_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_flush_iexec_1330_delayed_7_0_1249_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_flush_iexec_1330_delayed_7_0_1249_inst:started:   inputs: " & " flush_iexec_984 = "& Convert_SLV_To_Hex_String(flush_iexec_984));
          --
        end if; 
        if W_flush_iexec_1330_delayed_7_0_1249_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_flush_iexec_1330_delayed_7_0_1249_inst:finished:  outputs: " & " flush_iexec_1330_delayed_7_0_1251= "  & Convert_SLV_To_Hex_String(flush_iexec_1330_delayed_7_0_1251));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_flush_iexec_1330_delayed_7_0_1249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_flush_iexec_1330_delayed_7_0_1249_inst_req_0;
      W_flush_iexec_1330_delayed_7_0_1249_inst_ack_0<= wack(0);
      rreq(0) <= W_flush_iexec_1330_delayed_7_0_1249_inst_req_1;
      W_flush_iexec_1330_delayed_7_0_1249_inst_ack_1<= rack(0);
      W_flush_iexec_1330_delayed_7_0_1249_inst : InterlockBuffer generic map ( -- 
        name => "W_flush_iexec_1330_delayed_7_0_1249_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => flush_iexec_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => flush_iexec_1330_delayed_7_0_1251,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_icache_state_1063_delayed_7_0_1008_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_icache_state_1063_delayed_7_0_1008_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_icache_state_1063_delayed_7_0_1008_inst:started:   inputs: " & " icache_state_937 = "& Convert_SLV_To_Hex_String(icache_state_937));
          --
        end if; 
        if W_icache_state_1063_delayed_7_0_1008_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_icache_state_1063_delayed_7_0_1008_inst:finished:  outputs: " & " icache_state_1063_delayed_7_0_1010= "  & Convert_SLV_To_Hex_String(icache_state_1063_delayed_7_0_1010));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_icache_state_1063_delayed_7_0_1008_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_icache_state_1063_delayed_7_0_1008_inst_req_0;
      W_icache_state_1063_delayed_7_0_1008_inst_ack_0<= wack(0);
      rreq(0) <= W_icache_state_1063_delayed_7_0_1008_inst_req_1;
      W_icache_state_1063_delayed_7_0_1008_inst_ack_1<= rack(0);
      W_icache_state_1063_delayed_7_0_1008_inst : InterlockBuffer generic map ( -- 
        name => "W_icache_state_1063_delayed_7_0_1008_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 10,
        out_data_width => 10,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => icache_state_937,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => icache_state_1063_delayed_7_0_1010,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_idecode_state_1061_delayed_7_0_1005_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_idecode_state_1061_delayed_7_0_1005_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_idecode_state_1061_delayed_7_0_1005_inst:started:   inputs: " & " idecode_state_941 = "& Convert_SLV_To_Hex_String(idecode_state_941));
          --
        end if; 
        if W_idecode_state_1061_delayed_7_0_1005_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_idecode_state_1061_delayed_7_0_1005_inst:finished:  outputs: " & " idecode_state_1061_delayed_7_0_1007= "  & Convert_SLV_To_Hex_String(idecode_state_1061_delayed_7_0_1007));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_idecode_state_1061_delayed_7_0_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_idecode_state_1061_delayed_7_0_1005_inst_req_0;
      W_idecode_state_1061_delayed_7_0_1005_inst_ack_0<= wack(0);
      rreq(0) <= W_idecode_state_1061_delayed_7_0_1005_inst_req_1;
      W_idecode_state_1061_delayed_7_0_1005_inst_ack_1<= rack(0);
      W_idecode_state_1061_delayed_7_0_1005_inst : InterlockBuffer generic map ( -- 
        name => "W_idecode_state_1061_delayed_7_0_1005_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 42,
        out_data_width => 42,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => idecode_state_941,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idecode_state_1061_delayed_7_0_1007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iregfile_pc_1342_delayed_7_0_1261_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_iregfile_pc_1342_delayed_7_0_1261_inst:started:   inputs: " & " iregfile_pc_1034 = "& Convert_SLV_To_Hex_String(iregfile_pc_1034));
          --
        end if; 
        if W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_iregfile_pc_1342_delayed_7_0_1261_inst:finished:  outputs: " & " iregfile_pc_1342_delayed_7_0_1263= "  & Convert_SLV_To_Hex_String(iregfile_pc_1342_delayed_7_0_1263));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iregfile_pc_1342_delayed_7_0_1261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iregfile_pc_1342_delayed_7_0_1261_inst_req_0;
      W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_0<= wack(0);
      rreq(0) <= W_iregfile_pc_1342_delayed_7_0_1261_inst_req_1;
      W_iregfile_pc_1342_delayed_7_0_1261_inst_ack_1<= rack(0);
      W_iregfile_pc_1342_delayed_7_0_1261_inst : InterlockBuffer generic map ( -- 
        name => "W_iregfile_pc_1342_delayed_7_0_1261_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 10,
        out_data_width => 10,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iregfile_pc_1034,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iregfile_pc_1342_delayed_7_0_1263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst:started:   inputs: " & " iretire_state_to_rs1_imm_1191 = "& Convert_SLV_To_Hex_String(iretire_state_to_rs1_imm_1191));
          --
        end if; 
        if W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst:finished:  outputs: " & " iretire_state_to_rs1_imm_1318_delayed_7_0_1227= "  & Convert_SLV_To_Hex_String(iretire_state_to_rs1_imm_1318_delayed_7_0_1227));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_0;
      W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_0<= wack(0);
      rreq(0) <= W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_req_1;
      W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst_ack_1<= rack(0);
      W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst : InterlockBuffer generic map ( -- 
        name => "W_iretire_state_to_rs1_imm_1318_delayed_7_0_1225_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iretire_state_to_rs1_imm_1191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iretire_state_to_rs1_imm_1318_delayed_7_0_1227,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst:started:   inputs: " & " iretire_state_to_rs2_1195 = "& Convert_SLV_To_Hex_String(iretire_state_to_rs2_1195));
          --
        end if; 
        if W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst:finished:  outputs: " & " iretire_state_to_rs2_1324_delayed_7_0_1239= "  & Convert_SLV_To_Hex_String(iretire_state_to_rs2_1324_delayed_7_0_1239));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_0;
      W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_0<= wack(0);
      rreq(0) <= W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_req_1;
      W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst_ack_1<= rack(0);
      W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst : InterlockBuffer generic map ( -- 
        name => "W_iretire_state_to_rs2_1324_delayed_7_0_1237_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iretire_state_to_rs2_1195,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iretire_state_to_rs2_1324_delayed_7_0_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_reg_data_to_be_written_1212_inst flow-through 
    process(reg_data_to_be_written_1214) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_reg_data_to_be_written_1212_inst:flowthrough inputs: " & " iretire_exec_result_memData_1094 = "& Convert_SLV_To_Hex_String(iretire_exec_result_memData_1094) & " outputs:" & " reg_data_to_be_written_1214= "  & Convert_SLV_To_Hex_String(reg_data_to_be_written_1214));
      --
    end process; 
    -- interlock W_reg_data_to_be_written_1212_inst
    process(iretire_exec_result_memData_1094) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iretire_exec_result_memData_1094(31 downto 0);
      reg_data_to_be_written_1214 <= tmp_var; -- 
    end process;
    -- logger for split-operator W_reg_data_to_be_written_1319_delayed_7_0_1228_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_reg_data_to_be_written_1319_delayed_7_0_1228_inst:started:   inputs: " & " reg_data_to_be_written_1214 = "& Convert_SLV_To_Hex_String(reg_data_to_be_written_1214));
          --
        end if; 
        if W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_reg_data_to_be_written_1319_delayed_7_0_1228_inst:finished:  outputs: " & " reg_data_to_be_written_1319_delayed_7_0_1230= "  & Convert_SLV_To_Hex_String(reg_data_to_be_written_1319_delayed_7_0_1230));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_0;
      W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_0<= wack(0);
      rreq(0) <= W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_req_1;
      W_reg_data_to_be_written_1319_delayed_7_0_1228_inst_ack_1<= rack(0);
      W_reg_data_to_be_written_1319_delayed_7_0_1228_inst : InterlockBuffer generic map ( -- 
        name => "W_reg_data_to_be_written_1319_delayed_7_0_1228_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => reg_data_to_be_written_1214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => reg_data_to_be_written_1319_delayed_7_0_1230,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_reg_data_to_be_written_1325_delayed_7_0_1240_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_reg_data_to_be_written_1325_delayed_7_0_1240_inst:started:   inputs: " & " reg_data_to_be_written_1214 = "& Convert_SLV_To_Hex_String(reg_data_to_be_written_1214));
          --
        end if; 
        if W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_reg_data_to_be_written_1325_delayed_7_0_1240_inst:finished:  outputs: " & " reg_data_to_be_written_1325_delayed_7_0_1242= "  & Convert_SLV_To_Hex_String(reg_data_to_be_written_1325_delayed_7_0_1242));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_0;
      W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_0<= wack(0);
      rreq(0) <= W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_req_1;
      W_reg_data_to_be_written_1325_delayed_7_0_1240_inst_ack_1<= rack(0);
      W_reg_data_to_be_written_1325_delayed_7_0_1240_inst : InterlockBuffer generic map ( -- 
        name => "W_reg_data_to_be_written_1325_delayed_7_0_1240_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => reg_data_to_be_written_1214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => reg_data_to_be_written_1325_delayed_7_0_1242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_stall_first_4_1060_delayed_7_0_1002_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_stall_first_4_1060_delayed_7_0_1002_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_stall_first_4_1060_delayed_7_0_1002_inst:started:   inputs: " & " stall_first_4_984 = "& Convert_SLV_To_Hex_String(stall_first_4_984));
          --
        end if; 
        if W_stall_first_4_1060_delayed_7_0_1002_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:W_stall_first_4_1060_delayed_7_0_1002_inst:finished:  outputs: " & " stall_first_4_1060_delayed_7_0_1004= "  & Convert_SLV_To_Hex_String(stall_first_4_1060_delayed_7_0_1004));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_stall_first_4_1060_delayed_7_0_1002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_stall_first_4_1060_delayed_7_0_1002_inst_req_0;
      W_stall_first_4_1060_delayed_7_0_1002_inst_ack_0<= wack(0);
      rreq(0) <= W_stall_first_4_1060_delayed_7_0_1002_inst_req_1;
      W_stall_first_4_1060_delayed_7_0_1002_inst_ack_1<= rack(0);
      W_stall_first_4_1060_delayed_7_0_1002_inst : InterlockBuffer generic map ( -- 
        name => "W_stall_first_4_1060_delayed_7_0_1002_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => stall_first_4_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => stall_first_4_1060_delayed_7_0_1004,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_dcache_state_1142_956_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_dcache_state_1142_956_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_dcache_state_1142_956_buf:started:   inputs: " & " n_dcache_state_1142 = "& Convert_SLV_To_Hex_String(n_dcache_state_1142));
          --
        end if; 
        if n_dcache_state_1142_956_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_dcache_state_1142_956_buf:finished:  outputs: " & " n_dcache_state_1142_956_buffered= "  & Convert_SLV_To_Hex_String(n_dcache_state_1142_956_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_dcache_state_1142_956_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_dcache_state_1142_956_buf_req_0;
      n_dcache_state_1142_956_buf_ack_0<= wack(0);
      rreq(0) <= n_dcache_state_1142_956_buf_req_1;
      n_dcache_state_1142_956_buf_ack_1<= rack(0);
      n_dcache_state_1142_956_buf : InterlockBuffer generic map ( -- 
        name => "n_dcache_state_1142_956_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 139,
        out_data_width => 139,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_dcache_state_1142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_dcache_state_1142_956_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_iRetire_state_1317_960_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_iRetire_state_1317_960_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_iRetire_state_1317_960_buf:started:   inputs: " & " n_iRetire_state_1317 = "& Convert_SLV_To_Hex_String(n_iRetire_state_1317));
          --
        end if; 
        if n_iRetire_state_1317_960_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_iRetire_state_1317_960_buf:finished:  outputs: " & " n_iRetire_state_1317_960_buffered= "  & Convert_SLV_To_Hex_String(n_iRetire_state_1317_960_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_iRetire_state_1317_960_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_iRetire_state_1317_960_buf_req_0;
      n_iRetire_state_1317_960_buf_ack_0<= wack(0);
      rreq(0) <= n_iRetire_state_1317_960_buf_req_1;
      n_iRetire_state_1317_960_buf_ack_1<= rack(0);
      n_iRetire_state_1317_960_buf : InterlockBuffer generic map ( -- 
        name => "n_iRetire_state_1317_960_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 139,
        out_data_width => 139,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_iRetire_state_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_iRetire_state_1317_960_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_icache_state_998_940_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_icache_state_998_940_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_icache_state_998_940_buf:started:   inputs: " & " n_icache_state_998 = "& Convert_SLV_To_Hex_String(n_icache_state_998));
          --
        end if; 
        if n_icache_state_998_940_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_icache_state_998_940_buf:finished:  outputs: " & " n_icache_state_998_940_buffered= "  & Convert_SLV_To_Hex_String(n_icache_state_998_940_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_icache_state_998_940_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_icache_state_998_940_buf_req_0;
      n_icache_state_998_940_buf_ack_0<= wack(0);
      rreq(0) <= n_icache_state_998_940_buf_req_1;
      n_icache_state_998_940_buf_ack_1<= rack(0);
      n_icache_state_998_940_buf : InterlockBuffer generic map ( -- 
        name => "n_icache_state_998_940_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 10,
        out_data_width => 10,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_icache_state_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_icache_state_998_940_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_idecode_state_1021_944_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_idecode_state_1021_944_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_idecode_state_1021_944_buf:started:   inputs: " & " n_idecode_state_1021 = "& Convert_SLV_To_Hex_String(n_idecode_state_1021));
          --
        end if; 
        if n_idecode_state_1021_944_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_idecode_state_1021_944_buf:finished:  outputs: " & " n_idecode_state_1021_944_buffered= "  & Convert_SLV_To_Hex_String(n_idecode_state_1021_944_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_idecode_state_1021_944_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_idecode_state_1021_944_buf_req_0;
      n_idecode_state_1021_944_buf_ack_0<= wack(0);
      rreq(0) <= n_idecode_state_1021_944_buf_req_1;
      n_idecode_state_1021_944_buf_ack_1<= rack(0);
      n_idecode_state_1021_944_buf : InterlockBuffer generic map ( -- 
        name => "n_idecode_state_1021_944_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 42,
        out_data_width => 42,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_idecode_state_1021,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_idecode_state_1021_944_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_iexec_state_1275_952_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_iexec_state_1275_952_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_iexec_state_1275_952_buf:started:   inputs: " & " n_iexec_state_1275 = "& Convert_SLV_To_Hex_String(n_iexec_state_1275));
          --
        end if; 
        if n_iexec_state_1275_952_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_iexec_state_1275_952_buf:finished:  outputs: " & " n_iexec_state_1275_952_buffered= "  & Convert_SLV_To_Hex_String(n_iexec_state_1275_952_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_iexec_state_1275_952_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_iexec_state_1275_952_buf_req_0;
      n_iexec_state_1275_952_buf_ack_0<= wack(0);
      rreq(0) <= n_iexec_state_1275_952_buf_req_1;
      n_iexec_state_1275_952_buf_ack_1<= rack(0);
      n_iexec_state_1275_952_buf : InterlockBuffer generic map ( -- 
        name => "n_iexec_state_1275_952_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 106,
        out_data_width => 106,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_iexec_state_1275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_iexec_state_1275_952_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_iregfile_state_1030_948_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_iregfile_state_1030_948_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_iregfile_state_1030_948_buf:started:   inputs: " & " n_iregfile_state_1030 = "& Convert_SLV_To_Hex_String(n_iregfile_state_1030));
          --
        end if; 
        if n_iregfile_state_1030_948_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:n_iregfile_state_1030_948_buf:finished:  outputs: " & " n_iregfile_state_1030_948_buffered= "  & Convert_SLV_To_Hex_String(n_iregfile_state_1030_948_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_iregfile_state_1030_948_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_iregfile_state_1030_948_buf_req_0;
      n_iregfile_state_1030_948_buf_ack_0<= wack(0);
      rreq(0) <= n_iregfile_state_1030_948_buf_req_1;
      n_iregfile_state_1030_948_buf_ack_1<= rack(0);
      n_iregfile_state_1030_948_buf : InterlockBuffer generic map ( -- 
        name => "n_iregfile_state_1030_948_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 42,
        out_data_width => 42,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_iregfile_state_1030,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_iregfile_state_1030_948_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator next_ifetch_state_1358_936_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if next_ifetch_state_1358_936_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:next_ifetch_state_1358_936_buf:started:   inputs: " & " next_ifetch_state_1358 = "& Convert_SLV_To_Hex_String(next_ifetch_state_1358));
          --
        end if; 
        if next_ifetch_state_1358_936_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:next_ifetch_state_1358_936_buf:finished:  outputs: " & " next_ifetch_state_1358_936_buffered= "  & Convert_SLV_To_Hex_String(next_ifetch_state_1358_936_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    next_ifetch_state_1358_936_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_ifetch_state_1358_936_buf_req_0;
      next_ifetch_state_1358_936_buf_ack_0<= wack(0);
      rreq(0) <= next_ifetch_state_1358_936_buf_req_1;
      next_ifetch_state_1358_936_buf_ack_1<= rack(0);
      next_ifetch_state_1358_936_buf : InterlockBuffer generic map ( -- 
        name => "next_ifetch_state_1358_936_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 10,
        out_data_width => 10,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_ifetch_state_1358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_ifetch_state_1358_936_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1346_inst flow-through 
    process(type_cast_1346_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:type_cast_1346_inst:flowthrough inputs: " & " ifetch_state_933 = "& Convert_SLV_To_Hex_String(ifetch_state_933) & " outputs:" & " type_cast_1346_wire= "  & Convert_SLV_To_Hex_String(type_cast_1346_wire));
      --
    end process; 
    -- interlock type_cast_1346_inst
    process(ifetch_state_933) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 9 downto 0) := ifetch_state_933(9 downto 0);
      type_cast_1346_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1350_inst flow-through 
    process(type_cast_1350_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:type_cast_1350_inst:flowthrough inputs: " & " ADD_u10_u10_1349_wire = "& Convert_SLV_To_Hex_String(ADD_u10_u10_1349_wire) & " outputs:" & " type_cast_1350_wire= "  & Convert_SLV_To_Hex_String(type_cast_1350_wire));
      --
    end process; 
    -- interlock type_cast_1350_inst
    process(ADD_u10_u10_1349_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 9 downto 0) := ADD_u10_u10_1349_wire(9 downto 0);
      type_cast_1350_wire <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_931_branch_req_0," req0 do_while_stmt_931_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_931_branch_ack_0," ack0 do_while_stmt_931_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_931_branch_ack_1," ack1 do_while_stmt_931_branch");
    do_while_stmt_931_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1377_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_931_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_931_branch_req_0,
          ack0 => do_while_stmt_931_branch_ack_0,
          ack1 => do_while_stmt_931_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_926_branch_req_0," req0 if_stmt_926_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_926_branch_ack_0," ack0 if_stmt_926_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_926_branch_ack_1," ack1 if_stmt_926_branch");
    if_stmt_926_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u8_u1_929_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_926_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_926_branch_req_0,
          ack0 => if_stmt_926_branch_ack_0,
          ack1 => if_stmt_926_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u10_u10_1349_inst flow-through 
    process(ADD_u10_u10_1349_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:ADD_u10_u10_1349_inst:flowthrough inputs: " & " ifetch_state_933 = "& Convert_SLV_To_Hex_String(ifetch_state_933) & " konst_1348_wire_constant = "& Convert_SLV_To_Hex_String(konst_1348_wire_constant) & " outputs:" & " ADD_u10_u10_1349_wire= "  & Convert_SLV_To_Hex_String(ADD_u10_u10_1349_wire));
      --
    end process; 
    -- binary operator ADD_u10_u10_1349_inst
    process(ifetch_state_933) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ifetch_state_933, konst_1348_wire_constant, tmp_var);
      ADD_u10_u10_1349_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u24_1295_inst flow-through 
    process(CONCAT_u16_u24_1295_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u16_u24_1295_inst:flowthrough inputs: " & " CONCAT_u8_u16_1293_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_1293_wire) & " dcache_rs2_1058 = "& Convert_SLV_To_Hex_String(dcache_rs2_1058) & " outputs:" & " CONCAT_u16_u24_1295_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u24_1295_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u24_1295_inst
    process(CONCAT_u8_u16_1293_wire, dcache_rs2_1058) -- 
      variable tmp_var : std_logic_vector(23 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_1293_wire, dcache_rs2_1058, tmp_var);
      CONCAT_u16_u24_1295_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1259_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u16_u32_1259_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u16_u32_1259_inst:started:   inputs: " & " CONCAT_u8_u16_1255_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_1255_wire) & " CONCAT_u8_u16_1258_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_1258_wire));
          --
        end if; 
        if CONCAT_u16_u32_1259_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u16_u32_1259_inst:finished:  outputs: " & " CONCAT_u16_u32_1338_1338_delayed_7_0_1260= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1338_1338_delayed_7_0_1260));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (2) : CONCAT_u16_u32_1259_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_1255_wire & CONCAT_u8_u16_1258_wire;
      CONCAT_u16_u32_1338_1338_delayed_7_0_1260 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_1259_inst_req_0;
      CONCAT_u16_u32_1259_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_1259_inst_req_1;
      CONCAT_u16_u32_1259_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 7,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- logger for split-operator CONCAT_u1_u11_1307_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u1_u11_1307_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u1_u11_1307_inst:started:   inputs: " & " dcache_isBranch_1078 = "& Convert_SLV_To_Hex_String(dcache_isBranch_1078) & " dcache_pc_1082 = "& Convert_SLV_To_Hex_String(dcache_pc_1082));
          --
        end if; 
        if CONCAT_u1_u11_1307_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u1_u11_1307_inst:finished:  outputs: " & " CONCAT_u1_u11_1370_1370_delayed_7_0_1308= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u11_1370_1370_delayed_7_0_1308));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (3) : CONCAT_u1_u11_1307_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= dcache_isBranch_1078 & dcache_pc_1082;
      CONCAT_u1_u11_1370_1370_delayed_7_0_1308 <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u11_1307_inst_req_0;
      CONCAT_u1_u11_1307_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u11_1307_inst_req_1;
      CONCAT_u1_u11_1307_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 10, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 7,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- logger for split-operator CONCAT_u24_u64_1299_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u24_u64_1299_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u24_u64_1299_inst:started:   inputs: " & " CONCAT_u16_u24_1295_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u24_1295_wire) & " CONCAT_u8_u40_1298_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u40_1298_wire));
          --
        end if; 
        if CONCAT_u24_u64_1299_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u24_u64_1299_inst:finished:  outputs: " & " CONCAT_u24_u64_1364_1364_delayed_7_0_1300= "  & Convert_SLV_To_Hex_String(CONCAT_u24_u64_1364_1364_delayed_7_0_1300));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (4) : CONCAT_u24_u64_1299_inst 
    ApConcat_group_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u24_1295_wire & CONCAT_u8_u40_1298_wire;
      CONCAT_u24_u64_1364_1364_delayed_7_0_1300 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u24_u64_1299_inst_req_0;
      CONCAT_u24_u64_1299_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u24_u64_1299_inst_req_1;
      CONCAT_u24_u64_1299_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_4_gI: SplitGuardInterface generic map(name => "ApConcat_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 24,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 40, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 7,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- logger for split-operator CONCAT_u32_u106_1273_inst flow-through 
    process(CONCAT_u32_u106_1273_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u32_u106_1273_inst:flowthrough inputs: " & " CONCAT_u16_u32_1338_1338_delayed_7_0_1260 = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1338_1338_delayed_7_0_1260) & " CONCAT_u64_u74_1272_wire = "& Convert_SLV_To_Hex_String(CONCAT_u64_u74_1272_wire) & " outputs:" & " CONCAT_u32_u106_1273_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u106_1273_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u106_1273_inst
    process(CONCAT_u16_u32_1338_1338_delayed_7_0_1260, CONCAT_u64_u74_1272_wire) -- 
      variable tmp_var : std_logic_vector(105 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u32_1338_1338_delayed_7_0_1260, CONCAT_u64_u74_1272_wire, tmp_var);
      CONCAT_u32_u106_1273_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u42_1018_inst flow-through 
    process(CONCAT_u32_u42_1018_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u32_u42_1018_inst:flowthrough inputs: " & " icache_instruction_989 = "& Convert_SLV_To_Hex_String(icache_instruction_989) & " icache_state_1063_delayed_7_0_1010 = "& Convert_SLV_To_Hex_String(icache_state_1063_delayed_7_0_1010) & " outputs:" & " CONCAT_u32_u42_1018_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u42_1018_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u42_1018_inst
    process(icache_instruction_989, icache_state_1063_delayed_7_0_1010) -- 
      variable tmp_var : std_logic_vector(41 downto 0); -- 
    begin -- 
      ApConcat_proc(icache_instruction_989, icache_state_1063_delayed_7_0_1010, tmp_var);
      CONCAT_u32_u42_1018_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_1270_inst flow-through 
    process(CONCAT_u32_u64_1270_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u32_u64_1270_inst:flowthrough inputs: " & " final_rd1_1236 = "& Convert_SLV_To_Hex_String(final_rd1_1236) & " final_rd2_1248 = "& Convert_SLV_To_Hex_String(final_rd2_1248) & " outputs:" & " CONCAT_u32_u64_1270_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_1270_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_1270_inst
    process(final_rd1_1236, final_rd2_1248) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(final_rd1_1236, final_rd2_1248, tmp_var);
      CONCAT_u32_u64_1270_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_1313_inst flow-through 
    process(CONCAT_u32_u64_1313_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u32_u64_1313_inst:flowthrough inputs: " & " dcache_rd2_1365_delayed_7_0_1303 = "& Convert_SLV_To_Hex_String(dcache_rd2_1365_delayed_7_0_1303) & " dcache_data_to_be_written_to_reg_1289 = "& Convert_SLV_To_Hex_String(dcache_data_to_be_written_to_reg_1289) & " outputs:" & " CONCAT_u32_u64_1313_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_1313_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_1313_inst
    process(dcache_rd2_1365_delayed_7_0_1303, dcache_data_to_be_written_to_reg_1289) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(dcache_rd2_1365_delayed_7_0_1303, dcache_data_to_be_written_to_reg_1289, tmp_var);
      CONCAT_u32_u64_1313_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u64_u139_1316_inst flow-through 
    process(n_iRetire_state_1317) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u64_u139_1316_inst:flowthrough inputs: " & " CONCAT_u24_u64_1364_1364_delayed_7_0_1300 = "& Convert_SLV_To_Hex_String(CONCAT_u24_u64_1364_1364_delayed_7_0_1300) & " CONCAT_u64_u75_1315_wire = "& Convert_SLV_To_Hex_String(CONCAT_u64_u75_1315_wire) & " outputs:" & " n_iRetire_state_1317= "  & Convert_SLV_To_Hex_String(n_iRetire_state_1317));
      --
    end process; 
    -- binary operator CONCAT_u64_u139_1316_inst
    process(CONCAT_u24_u64_1364_1364_delayed_7_0_1300, CONCAT_u64_u75_1315_wire) -- 
      variable tmp_var : std_logic_vector(138 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u24_u64_1364_1364_delayed_7_0_1300, CONCAT_u64_u75_1315_wire, tmp_var);
      n_iRetire_state_1317 <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u64_u74_1272_inst flow-through 
    process(CONCAT_u64_u74_1272_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u64_u74_1272_inst:flowthrough inputs: " & " CONCAT_u32_u64_1270_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_1270_wire) & " iregfile_pc_1342_delayed_7_0_1263 = "& Convert_SLV_To_Hex_String(iregfile_pc_1342_delayed_7_0_1263) & " outputs:" & " CONCAT_u64_u74_1272_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u64_u74_1272_wire));
      --
    end process; 
    -- binary operator CONCAT_u64_u74_1272_inst
    process(CONCAT_u32_u64_1270_wire, iregfile_pc_1342_delayed_7_0_1263) -- 
      variable tmp_var : std_logic_vector(73 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_1270_wire, iregfile_pc_1342_delayed_7_0_1263, tmp_var);
      CONCAT_u64_u74_1272_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u64_u75_1315_inst flow-through 
    process(CONCAT_u64_u75_1315_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u64_u75_1315_inst:flowthrough inputs: " & " CONCAT_u32_u64_1313_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_1313_wire) & " CONCAT_u1_u11_1370_1370_delayed_7_0_1308 = "& Convert_SLV_To_Hex_String(CONCAT_u1_u11_1370_1370_delayed_7_0_1308) & " outputs:" & " CONCAT_u64_u75_1315_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u64_u75_1315_wire));
      --
    end process; 
    -- binary operator CONCAT_u64_u75_1315_inst
    process(CONCAT_u32_u64_1313_wire, CONCAT_u1_u11_1370_1370_delayed_7_0_1308) -- 
      variable tmp_var : std_logic_vector(74 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_1313_wire, CONCAT_u1_u11_1370_1370_delayed_7_0_1308, tmp_var);
      CONCAT_u64_u75_1315_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u8_u16_1255_inst flow-through 
    process(CONCAT_u8_u16_1255_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u8_u16_1255_inst:flowthrough inputs: " & " reg_opcode_1199 = "& Convert_SLV_To_Hex_String(reg_opcode_1199) & " reg_rs1_imm_1203 = "& Convert_SLV_To_Hex_String(reg_rs1_imm_1203) & " outputs:" & " CONCAT_u8_u16_1255_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_1255_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_1255_inst
    process(reg_opcode_1199, reg_rs1_imm_1203) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(reg_opcode_1199, reg_rs1_imm_1203, tmp_var);
      CONCAT_u8_u16_1255_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u8_u16_1258_inst flow-through 
    process(CONCAT_u8_u16_1258_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u8_u16_1258_inst:flowthrough inputs: " & " reg_rs2_1207 = "& Convert_SLV_To_Hex_String(reg_rs2_1207) & " reg_rd_1211 = "& Convert_SLV_To_Hex_String(reg_rd_1211) & " outputs:" & " CONCAT_u8_u16_1258_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_1258_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_1258_inst
    process(reg_rs2_1207, reg_rd_1211) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(reg_rs2_1207, reg_rd_1211, tmp_var);
      CONCAT_u8_u16_1258_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u8_u16_1293_inst flow-through 
    process(CONCAT_u8_u16_1293_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u8_u16_1293_inst:flowthrough inputs: " & " dcache_opcode_1050 = "& Convert_SLV_To_Hex_String(dcache_opcode_1050) & " dcache_rs1_imm_1054 = "& Convert_SLV_To_Hex_String(dcache_rs1_imm_1054) & " outputs:" & " CONCAT_u8_u16_1293_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_1293_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_1293_inst
    process(dcache_opcode_1050, dcache_rs1_imm_1054) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(dcache_opcode_1050, dcache_rs1_imm_1054, tmp_var);
      CONCAT_u8_u16_1293_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u8_u40_1298_inst flow-through 
    process(CONCAT_u8_u40_1298_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:CONCAT_u8_u40_1298_inst:flowthrough inputs: " & " dcache_rd_1062 = "& Convert_SLV_To_Hex_String(dcache_rd_1062) & " dcache_rd1_1066 = "& Convert_SLV_To_Hex_String(dcache_rd1_1066) & " outputs:" & " CONCAT_u8_u40_1298_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u40_1298_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u40_1298_inst
    process(dcache_rd_1062, dcache_rd1_1066) -- 
      variable tmp_var : std_logic_vector(39 downto 0); -- 
    begin -- 
      ApConcat_proc(dcache_rd_1062, dcache_rd1_1066, tmp_var);
      CONCAT_u8_u40_1298_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_1279_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if EQ_u8_u1_1279_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:EQ_u8_u1_1279_inst:started:   inputs: " & " dcache_opcode_1050 = "& Convert_SLV_To_Hex_String(dcache_opcode_1050) & " R_LOAD_1278_wire_constant = "& Convert_SLV_To_Hex_String(R_LOAD_1278_wire_constant));
          --
        end if; 
        if EQ_u8_u1_1279_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:EQ_u8_u1_1279_inst:finished:  outputs: " & " EQ_u8_u1_1350_1350_delayed_7_0_1280= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_1350_1350_delayed_7_0_1280));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (16) : EQ_u8_u1_1279_inst 
    ApIntEq_group_16: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= dcache_opcode_1050;
      EQ_u8_u1_1350_1350_delayed_7_0_1280 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_1279_inst_req_0;
      EQ_u8_u1_1279_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_1279_inst_req_1;
      EQ_u8_u1_1279_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_16_gI: SplitGuardInterface generic map(name => "ApIntEq_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          buffering  => 7,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- logger for split-operator EQ_u8_u1_1321_inst flow-through 
    process(EQ_u8_u1_1321_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:EQ_u8_u1_1321_inst:flowthrough inputs: " & " dcache_rs2_1058 = "& Convert_SLV_To_Hex_String(dcache_rs2_1058) & " iretire_rd_1090 = "& Convert_SLV_To_Hex_String(iretire_rd_1090) & " outputs:" & " EQ_u8_u1_1321_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_1321_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_1321_inst
    process(dcache_rs2_1058, iretire_rd_1090) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_rs2_1058, iretire_rd_1090, tmp_var);
      EQ_u8_u1_1321_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_1329_inst flow-through 
    process(EQ_u8_u1_1329_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:EQ_u8_u1_1329_inst:flowthrough inputs: " & " dcache_rd_1062 = "& Convert_SLV_To_Hex_String(dcache_rd_1062) & " iexec_rs1_imm_1038 = "& Convert_SLV_To_Hex_String(iexec_rs1_imm_1038) & " outputs:" & " EQ_u8_u1_1329_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_1329_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_1329_inst
    process(dcache_rd_1062, iexec_rs1_imm_1038) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_rd_1062, iexec_rs1_imm_1038, tmp_var);
      EQ_u8_u1_1329_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_1333_inst flow-through 
    process(EQ_u8_u1_1333_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:EQ_u8_u1_1333_inst:flowthrough inputs: " & " iretire_rd_1090 = "& Convert_SLV_To_Hex_String(iretire_rd_1090) & " iexec_rs1_imm_1038 = "& Convert_SLV_To_Hex_String(iexec_rs1_imm_1038) & " outputs:" & " EQ_u8_u1_1333_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_1333_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_1333_inst
    process(iretire_rd_1090, iexec_rs1_imm_1038) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_rd_1090, iexec_rs1_imm_1038, tmp_var);
      EQ_u8_u1_1333_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_1376_inst flow-through 
    process(EQ_u8_u1_1376_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:EQ_u8_u1_1376_inst:flowthrough inputs: " & " iretire_opcode_1086 = "& Convert_SLV_To_Hex_String(iretire_opcode_1086) & " R_HALT_1375_wire_constant = "& Convert_SLV_To_Hex_String(R_HALT_1375_wire_constant) & " outputs:" & " EQ_u8_u1_1376_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_1376_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_1376_inst
    process(iretire_opcode_1086) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_1086, R_HALT_1375_wire_constant, tmp_var);
      EQ_u8_u1_1376_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_929_inst flow-through 
    process(EQ_u8_u1_929_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:EQ_u8_u1_929_inst:flowthrough inputs: " & " cmd_925 = "& Convert_SLV_To_Hex_String(cmd_925) & " R_one_8_928_wire_constant = "& Convert_SLV_To_Hex_String(R_one_8_928_wire_constant) & " outputs:" & " EQ_u8_u1_929_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_929_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_929_inst
    process(cmd_925) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(cmd_925, R_one_8_928_wire_constant, tmp_var);
      EQ_u8_u1_929_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_1377_inst flow-through 
    process(NOT_u1_u1_1377_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:NOT_u1_u1_1377_inst:flowthrough inputs: " & " EQ_u8_u1_1376_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_1376_wire) & " outputs:" & " NOT_u1_u1_1377_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_1377_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_1377_inst
    process(EQ_u8_u1_1376_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", EQ_u8_u1_1376_wire, tmp_var);
      NOT_u1_u1_1377_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator RPIPE_start_processor_924_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_start_processor_924_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:RPIPE_start_processor_924_inst:started:   PipeRead from start_processor inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_start_processor_924_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:RPIPE_start_processor_924_inst:finished:  outputs: " & " cmd_925= "  & Convert_SLV_To_Hex_String(cmd_925));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_start_processor_924_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_start_processor_924_inst_req_0;
      RPIPE_start_processor_924_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_start_processor_924_inst_req_1;
      RPIPE_start_processor_924_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      cmd_925 <= data_out(7 downto 0);
      start_processor_read_0_gI: SplitGuardInterface generic map(name => "start_processor_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      start_processor_read_0: InputPortRevised -- 
        generic map ( name => "start_processor_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => start_processor_pipe_read_req(0),
          oack => start_processor_pipe_read_ack(0),
          odata => start_processor_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_processor_result_1370_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_processor_result_1370_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:WPIPE_processor_result_1370_inst:started:   PipeWrite to processor_result inputs: " & " reg_data_to_be_written_1214 = "& Convert_SLV_To_Hex_String(reg_data_to_be_written_1214));
          --
        end if; 
        if WPIPE_processor_result_1370_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:WPIPE_processor_result_1370_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_processor_result_1370_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_processor_result_1370_inst_req_0;
      WPIPE_processor_result_1370_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_processor_result_1370_inst_req_1;
      WPIPE_processor_result_1370_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= reg_data_to_be_written_1214;
      processor_result_write_0_gI: SplitGuardInterface generic map(name => "processor_result_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      processor_result_write_0: OutputPortRevised -- 
        generic map ( name => "processor_result", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => processor_result_pipe_write_req(0),
          oack => processor_result_pipe_write_ack(0),
          odata => processor_result_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_1133_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1133_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_1133_call:started:  Call to module iExecStage inputs: " & " iexec_state_949 = "& Convert_SLV_To_Hex_String(iexec_state_949) & " iexec_rd1_final_1119 = "& Convert_SLV_To_Hex_String(iexec_rd1_final_1119) & " iexec_rd2_final_1128 = "& Convert_SLV_To_Hex_String(iexec_rd2_final_1128));
          --
        end if; 
        if call_stmt_1133_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_1133_call:finished:  outputs: " & " n_dcache_state_from_exec_1133= "  & Convert_SLV_To_Hex_String(n_dcache_state_from_exec_1133));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1133_call 
    iExecStage_call_group_0: Block -- 
      signal data_in: std_logic_vector(169 downto 0);
      signal data_out: std_logic_vector(138 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1133_call_req_0;
      call_stmt_1133_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1133_call_req_1;
      call_stmt_1133_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      iExecStage_call_group_0_gI: SplitGuardInterface generic map(name => "iExecStage_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iexec_state_949 & iexec_rd1_final_1119 & iexec_rd2_final_1128;
      n_dcache_state_from_exec_1133 <= data_out(138 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 170,
        owidth => 170,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => iExecStage_call_reqs(0),
          ackR => iExecStage_call_acks(0),
          dataR => iExecStage_call_data(169 downto 0),
          tagR => iExecStage_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 139,
          owidth => 139,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => iExecStage_return_acks(0), -- cross-over
          ackL => iExecStage_return_reqs(0), -- cross-over
          dataL => iExecStage_return_data(138 downto 0),
          tagL => iExecStage_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_989_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_989_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_989_call:started:  Call to module accessMem inputs: " & " R_read_signal_985_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_985_wire_constant) & " icache_state_937 = "& Convert_SLV_To_Hex_String(icache_state_937) & " R_zero_32_987_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_32_987_wire_constant));
          --
        end if; 
        if call_stmt_989_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_989_call:finished:  outputs: " & " icache_instruction_989= "  & Convert_SLV_To_Hex_String(icache_instruction_989));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_1175_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1175_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_1175_call:started:  Call to module accessMem inputs: " & " memWrite_1146 = "& Convert_SLV_To_Hex_String(memWrite_1146) & " memAddr_1170 = "& Convert_SLV_To_Hex_String(memAddr_1170) & " memWriteData_1160 = "& Convert_SLV_To_Hex_String(memWriteData_1160));
          --
        end if; 
        if call_stmt_1175_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_1175_call:finished:  outputs: " & " memReadData_1175= "  & Convert_SLV_To_Hex_String(memReadData_1175));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_989_call call_stmt_1175_call 
    accessMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 7, 1 => 7);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_989_call_req_0;
      reqL_unguarded(0) <= call_stmt_1175_call_req_0;
      call_stmt_989_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1175_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_989_call_req_1;
      reqR_unguarded(0) <= call_stmt_1175_call_req_1;
      call_stmt_989_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1175_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMem_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "accessMem_call_group_1_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMem_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "accessMem_call_group_1_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMem_call_group_1_gI: SplitGuardInterface generic map(name => "accessMem_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_read_signal_985_wire_constant & icache_state_937 & R_zero_32_987_wire_constant & memWrite_1146 & memAddr_1170 & memWriteData_1160;
      icache_instruction_989 <= data_out(63 downto 32);
      memReadData_1175 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(42 downto 0),
          tagR => accessMem_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(31 downto 0),
          tagL => accessMem_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_1224_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1224_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_1224_call:started:  Call to module accessReg inputs: " & " reg_valid_read1_1179 = "& Convert_SLV_To_Hex_String(reg_valid_read1_1179) & " reg_rs1_imm_1203 = "& Convert_SLV_To_Hex_String(reg_rs1_imm_1203) & " reg_valid_read2_1183 = "& Convert_SLV_To_Hex_String(reg_valid_read2_1183) & " reg_rs2_1207 = "& Convert_SLV_To_Hex_String(reg_rs2_1207) & " reg_valid_write_1187 = "& Convert_SLV_To_Hex_String(reg_valid_write_1187) & " iretire_rd_1090 = "& Convert_SLV_To_Hex_String(iretire_rd_1090) & " reg_data_to_be_written_1214 = "& Convert_SLV_To_Hex_String(reg_data_to_be_written_1214));
          --
        end if; 
        if call_stmt_1224_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_1224_call:finished:  outputs: " & " reg_d1_1224= "  & Convert_SLV_To_Hex_String(reg_d1_1224) & " reg_d2_1224= "  & Convert_SLV_To_Hex_String(reg_d2_1224));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_1224_call 
    accessReg_call_group_2: Block -- 
      signal data_in: std_logic_vector(58 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 7);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1224_call_req_0;
      call_stmt_1224_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1224_call_req_1;
      call_stmt_1224_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessReg_call_group_2_gI: SplitGuardInterface generic map(name => "accessReg_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= reg_valid_read1_1179 & reg_rs1_imm_1203 & reg_valid_read2_1183 & reg_rs2_1207 & reg_valid_write_1187 & iretire_rd_1090 & reg_data_to_be_written_1214;
      reg_d1_1224 <= data_out(63 downto 32);
      reg_d2_1224 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 59,
        owidth => 59,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessReg_call_reqs(0),
          ackR => accessReg_call_acks(0),
          dataR => accessReg_call_data(58 downto 0),
          tagR => accessReg_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessReg_return_acks(0), -- cross-over
          ackL => accessReg_return_reqs(0), -- cross-over
          dataL => accessReg_return_data(63 downto 0),
          tagL => accessReg_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- logger for split-operator call_stmt_984_call flow-through 
    process(ifetch_actions_984, icache_actions_984, idecode_actions_984, iregfile_actions_984, iexec_actions_984, dcache_actions_984, ex_Unconditional_JUMP_984, is_Branch_Hazard_984, flush_ifetch_984, flush_icache_984, flush_idecode_984, flush_reg_984, flush_iexec_984, flush_dcache_984, stall_first_4_984) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processor_daemon:DP:call_stmt_984_call:flowthrough inputs: " & " ifetch_state_933 = "& Convert_SLV_To_Hex_String(ifetch_state_933) & " icache_state_937 = "& Convert_SLV_To_Hex_String(icache_state_937) & " idecode_state_941 = "& Convert_SLV_To_Hex_String(idecode_state_941) & " iregfile_state_945 = "& Convert_SLV_To_Hex_String(iregfile_state_945) & " iexec_state_949 = "& Convert_SLV_To_Hex_String(iexec_state_949) & " dcache_state_953 = "& Convert_SLV_To_Hex_String(dcache_state_953) & " iretire_state_957 = "& Convert_SLV_To_Hex_String(iretire_state_957) & " outputs:" & " ifetch_actions_984= "  & Convert_SLV_To_Hex_String(ifetch_actions_984) & " icache_actions_984= "  & Convert_SLV_To_Hex_String(icache_actions_984) & " idecode_actions_984= "  & Convert_SLV_To_Hex_String(idecode_actions_984) & " iregfile_actions_984= "  & Convert_SLV_To_Hex_String(iregfile_actions_984) & " iexec_actions_984= "  & Convert_SLV_To_Hex_String(iexec_actions_984) & " dcache_actions_984= "  & Convert_SLV_To_Hex_String(dcache_actions_984) & " ex_Unconditional_JUMP_984= "  & Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_984) & " is_Branch_Hazard_984= "  & Convert_SLV_To_Hex_String(is_Branch_Hazard_984) & " flush_ifetch_984= "  & Convert_SLV_To_Hex_String(flush_ifetch_984) & " flush_icache_984= "  & Convert_SLV_To_Hex_String(flush_icache_984) & " flush_idecode_984= "  & Convert_SLV_To_Hex_String(flush_idecode_984) & " flush_reg_984= "  & Convert_SLV_To_Hex_String(flush_reg_984) & " flush_iexec_984= "  & Convert_SLV_To_Hex_String(flush_iexec_984) & " flush_dcache_984= "  & Convert_SLV_To_Hex_String(flush_dcache_984) & " stall_first_4_984= "  & Convert_SLV_To_Hex_String(stall_first_4_984));
      --
    end process; 
    volatile_operator_scoreBoard_2756: scoreBoard_Volatile port map(ifetch_state => ifetch_state_933, icache_state => icache_state_937, idecode_state => idecode_state_941, iregfile_state => iregfile_state_945, iexec_state => iexec_state_949, dcache_state => dcache_state_953, iretire_state => iretire_state_957, ifetch_actions => ifetch_actions_984, icache_actions => icache_actions_984, idecode_actions => idecode_actions_984, iregfile_actions => iregfile_actions_984, iexec_actions => iexec_actions_984, dcache_actions => dcache_actions_984, ex_Unconditional_JUMP => ex_Unconditional_JUMP_984, is_Branch_Hazard => is_Branch_Hazard_984, flush_ifetch => flush_ifetch_984, flush_icache => flush_icache_984, flush_idecode => flush_idecode_984, flush_reg => flush_reg_984, flush_iexec => flush_iexec_984, flush_dcache => flush_dcache_984, stall_first_4 => stall_first_4_984, clk => clk, reset => reset); 
    -- 
  end Block; -- data_path
  -- 
end processor_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity regAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    accessReg_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    accessReg_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    accessReg_request_pipe_read_data : in   std_logic_vector(63 downto 0);
    accessReg_response1_pipe_write_req : out  std_logic_vector(0 downto 0);
    accessReg_response1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    accessReg_response1_pipe_write_data : out  std_logic_vector(31 downto 0);
    accessReg_response2_pipe_write_req : out  std_logic_vector(0 downto 0);
    accessReg_response2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    accessReg_response2_pipe_write_data : out  std_logic_vector(31 downto 0);
    accessReg_call_reqs : out  std_logic_vector(0 downto 0);
    accessReg_call_acks : in   std_logic_vector(0 downto 0);
    accessReg_call_data : out  std_logic_vector(58 downto 0);
    accessReg_call_tag  :  out  std_logic_vector(0 downto 0);
    accessReg_return_reqs : out  std_logic_vector(0 downto 0);
    accessReg_return_acks : in   std_logic_vector(0 downto 0);
    accessReg_return_data : in   std_logic_vector(63 downto 0);
    accessReg_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity regAccessDaemon;
architecture regAccessDaemon_arch of regAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal regAccessDaemon_CP_1645_start: Boolean;
  signal regAccessDaemon_CP_1645_symbol: Boolean;
  -- volatile/operator module components. 
  component accessReg is -- 
    generic (tag_length : integer); 
    port ( -- 
      valid_1 : in  std_logic_vector(0 downto 0);
      addr_1 : in  std_logic_vector(7 downto 0);
      valid_2 : in  std_logic_vector(0 downto 0);
      addr_2 : in  std_logic_vector(7 downto 0);
      valid_w : in  std_logic_vector(0 downto 0);
      addr_w : in  std_logic_vector(7 downto 0);
      data_to_be_written : in  std_logic_vector(31 downto 0);
      read_data_1 : out  std_logic_vector(31 downto 0);
      read_data_2 : out  std_logic_vector(31 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1427_call_req_1 : boolean;
  signal call_stmt_1427_call_ack_1 : boolean;
  signal call_stmt_1427_call_req_0 : boolean;
  signal call_stmt_1427_call_ack_0 : boolean;
  signal RPIPE_accessReg_request_1388_inst_ack_1 : boolean;
  signal RPIPE_accessReg_request_1388_inst_req_1 : boolean;
  signal RPIPE_accessReg_request_1388_inst_ack_0 : boolean;
  signal RPIPE_accessReg_request_1388_inst_req_0 : boolean;
  signal do_while_stmt_1385_branch_req_0 : boolean;
  signal WPIPE_accessReg_response1_1428_inst_req_0 : boolean;
  signal WPIPE_accessReg_response1_1428_inst_ack_0 : boolean;
  signal WPIPE_accessReg_response1_1428_inst_req_1 : boolean;
  signal WPIPE_accessReg_response1_1428_inst_ack_1 : boolean;
  signal WPIPE_accessReg_response2_1431_inst_req_0 : boolean;
  signal WPIPE_accessReg_response2_1431_inst_ack_0 : boolean;
  signal WPIPE_accessReg_response2_1431_inst_req_1 : boolean;
  signal WPIPE_accessReg_response2_1431_inst_ack_1 : boolean;
  signal do_while_stmt_1385_branch_ack_0 : boolean;
  signal do_while_stmt_1385_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "regAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  regAccessDaemon_CP_1645_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "regAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= regAccessDaemon_CP_1645_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= regAccessDaemon_CP_1645_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= regAccessDaemon_CP_1645_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,regAccessDaemon_CP_1645_start,"regAccessDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,regAccessDaemon_CP_1645_symbol, "regAccessDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  regAccessDaemon_CP_1645: Block -- control-path 
    signal regAccessDaemon_CP_1645_elements: BooleanArray(28 downto 0);
    -- 
  begin -- 
    regAccessDaemon_CP_1645_elements(0) <= regAccessDaemon_CP_1645_start;
    regAccessDaemon_CP_1645_symbol <= regAccessDaemon_CP_1645_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1384/do_while_stmt_1385__entry__
      -- CP-element group 0: 	 branch_block_stmt_1384/branch_block_stmt_1384__entry__
      -- CP-element group 0: 	 branch_block_stmt_1384/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	28 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1384/do_while_stmt_1385__exit__
      -- CP-element group 1: 	 branch_block_stmt_1384/branch_block_stmt_1384__exit__
      -- CP-element group 1: 	 branch_block_stmt_1384/$exit
      -- CP-element group 1: 	 $exit
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_CP_1645_elements(1) <= regAccessDaemon_CP_1645_elements(28);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385__entry__
      -- CP-element group 2: 	 branch_block_stmt_1384/do_while_stmt_1385/$entry
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_CP_1645_elements(2) <= regAccessDaemon_CP_1645_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	28 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385__exit__
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group regAccessDaemon_CP_1645_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_back
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group regAccessDaemon_CP_1645_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	24 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	26 
    -- CP-element group 5: 	27 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1384/do_while_stmt_1385/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_taken/$entry
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_CP_1645_elements(5) <= regAccessDaemon_CP_1645_elements(24);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	25 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_body_done
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_CP_1645_elements(6) <= regAccessDaemon_CP_1645_elements(25);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_CP_1645_elements(7) <= regAccessDaemon_CP_1645_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_CP_1645_elements(8) <= regAccessDaemon_CP_1645_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	24 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/loop_body_start
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group regAccessDaemon_CP_1645_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_sample_start_
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:RPIPE_accessReg_request_1388_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(10), ack => RPIPE_accessReg_request_1388_inst_req_0); -- 
    regAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "regAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= regAccessDaemon_CP_1645_elements(9) & regAccessDaemon_CP_1645_elements(13);
      gj_regAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_update_start_
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:RPIPE_accessReg_request_1388_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(11), ack => RPIPE_accessReg_request_1388_inst_req_1); -- 
    regAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "regAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= regAccessDaemon_CP_1645_elements(12) & regAccessDaemon_CP_1645_elements(16);
      gj_regAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_sample_completed_
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:RPIPE_accessReg_request_1388_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_accessReg_request_1388_inst_ack_0, ack => regAccessDaemon_CP_1645_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/RPIPE_accessReg_request_1388_update_completed_
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:RPIPE_accessReg_request_1388_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_accessReg_request_1388_inst_ack_1, ack => regAccessDaemon_CP_1645_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Sample/crr
      -- CP-element group 14: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Sample/$entry
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:call_stmt_1427_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(14), ack => call_stmt_1427_call_req_0); -- 
    regAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "regAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= regAccessDaemon_CP_1645_elements(13) & regAccessDaemon_CP_1645_elements(16);
      gj_regAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	22 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Update/ccr
      -- CP-element group 15: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_update_start_
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:call_stmt_1427_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(15), ack => call_stmt_1427_call_req_1); -- 
    regAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "regAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= regAccessDaemon_CP_1645_elements(19) & regAccessDaemon_CP_1645_elements(22);
      gj_regAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Sample/cra
      -- CP-element group 16: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_sample_completed_
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:call_stmt_1427_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1427_call_ack_0, ack => regAccessDaemon_CP_1645_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_Update/cca
      -- CP-element group 17: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/call_stmt_1427_update_completed_
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:call_stmt_1427_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1427_call_ack_1, ack => regAccessDaemon_CP_1645_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Sample/req
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response1_1428_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(18), ack => WPIPE_accessReg_response1_1428_inst_req_0); -- 
    regAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "regAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= regAccessDaemon_CP_1645_elements(17) & regAccessDaemon_CP_1645_elements(20);
      gj_regAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Sample/ack
      -- CP-element group 19: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Update/req
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response1_1428_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response1_1428_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accessReg_response1_1428_inst_ack_0, ack => regAccessDaemon_CP_1645_elements(19)); -- 
    req_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(19), ack => WPIPE_accessReg_response1_1428_inst_req_1); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	25 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response1_1428_Update/ack
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response1_1428_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accessReg_response1_1428_inst_ack_1, ack => regAccessDaemon_CP_1645_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Sample/req
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response2_1431_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(21), ack => WPIPE_accessReg_response2_1431_inst_req_0); -- 
    regAccessDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "regAccessDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= regAccessDaemon_CP_1645_elements(17) & regAccessDaemon_CP_1645_elements(23);
      gj_regAccessDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	15 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Sample/ack
      -- CP-element group 22: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Update/req
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response2_1431_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response2_1431_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accessReg_response2_1431_inst_ack_0, ack => regAccessDaemon_CP_1645_elements(22)); -- 
    req_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(22), ack => WPIPE_accessReg_response2_1431_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/WPIPE_accessReg_response2_1431_Update/ack
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:WPIPE_accessReg_response2_1431_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accessReg_response2_1431_inst_ack_1, ack => regAccessDaemon_CP_1645_elements(23)); -- 
    -- CP-element group 24:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	9 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	5 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/condition_evaluated
      -- CP-element group 24: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:do_while_stmt_1385_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => regAccessDaemon_CP_1645_elements(24), ack => do_while_stmt_1385_branch_req_0); -- 
    -- Element group regAccessDaemon_CP_1645_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => regAccessDaemon_CP_1645_elements(9), ack => regAccessDaemon_CP_1645_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	6 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1384/do_while_stmt_1385/do_while_stmt_1385_loop_body/$exit
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 20);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "regAccessDaemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= regAccessDaemon_CP_1645_elements(20) & regAccessDaemon_CP_1645_elements(23);
      gj_regAccessDaemon_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	5 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_exit/$exit
      -- CP-element group 26: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_exit/ack
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:do_while_stmt_1385_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1385_branch_ack_0, ack => regAccessDaemon_CP_1645_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	5 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_taken/$exit
      -- CP-element group 27: 	 branch_block_stmt_1384/do_while_stmt_1385/loop_taken/ack
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:do_while_stmt_1385_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1385_branch_ack_1, ack => regAccessDaemon_CP_1645_elements(27)); -- 
    -- CP-element group 28:  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	3 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	1 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1384/do_while_stmt_1385/$exit
      -- 
    -- logger for CP element group regAccessDaemon_CP_1645_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and regAccessDaemon_CP_1645_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:regAccessDaemon:CP:regAccessDaemon_CP_1645_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    regAccessDaemon_CP_1645_elements(28) <= regAccessDaemon_CP_1645_elements(3);
    regAccessDaemon_do_while_stmt_1385_terminator_1736: loop_terminator -- 
      generic map (name => " regAccessDaemon_do_while_stmt_1385_terminator_1736", max_iterations_in_flight =>20) 
      port map(loop_body_exit => regAccessDaemon_CP_1645_elements(6),loop_continue => regAccessDaemon_CP_1645_elements(27),loop_terminate => regAccessDaemon_CP_1645_elements(26),loop_back => regAccessDaemon_CP_1645_elements(4),loop_exit => regAccessDaemon_CP_1645_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_1670_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= regAccessDaemon_CP_1645_elements(7);
        preds(1)  <= regAccessDaemon_CP_1645_elements(8);
        entry_tmerge_1670 : transition_merge -- 
          generic map(name => " entry_tmerge_1670")
          port map (preds => preds, symbol_out => regAccessDaemon_CP_1645_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addr1_1397 : std_logic_vector(7 downto 0);
    signal addr2_1405 : std_logic_vector(7 downto 0);
    signal addr_w_1413 : std_logic_vector(7 downto 0);
    signal cmd_1_1389 : std_logic_vector(63 downto 0);
    signal data_to_be_written_1417 : std_logic_vector(31 downto 0);
    signal konst_1435_wire_constant : std_logic_vector(0 downto 0);
    signal rdata1_1427 : std_logic_vector(31 downto 0);
    signal rdata2_1427 : std_logic_vector(31 downto 0);
    signal valid_1_1393 : std_logic_vector(0 downto 0);
    signal valid_2_1401 : std_logic_vector(0 downto 0);
    signal valid_w_1409 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1435_wire_constant <= "1";
    -- logger for split-operator slice_1392_inst flow-through 
    process(valid_1_1393) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:slice_1392_inst:flowthrough inputs: " & " cmd_1_1389 = "& Convert_SLV_To_Hex_String(cmd_1_1389) & " outputs:" & " valid_1_1393= "  & Convert_SLV_To_Hex_String(valid_1_1393));
      --
    end process; 
    -- flow-through slice operator slice_1392_inst
    valid_1_1393 <= cmd_1_1389(63 downto 63);
    -- logger for split-operator slice_1396_inst flow-through 
    process(addr1_1397) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:slice_1396_inst:flowthrough inputs: " & " cmd_1_1389 = "& Convert_SLV_To_Hex_String(cmd_1_1389) & " outputs:" & " addr1_1397= "  & Convert_SLV_To_Hex_String(addr1_1397));
      --
    end process; 
    -- flow-through slice operator slice_1396_inst
    addr1_1397 <= cmd_1_1389(62 downto 55);
    -- logger for split-operator slice_1400_inst flow-through 
    process(valid_2_1401) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:slice_1400_inst:flowthrough inputs: " & " cmd_1_1389 = "& Convert_SLV_To_Hex_String(cmd_1_1389) & " outputs:" & " valid_2_1401= "  & Convert_SLV_To_Hex_String(valid_2_1401));
      --
    end process; 
    -- flow-through slice operator slice_1400_inst
    valid_2_1401 <= cmd_1_1389(54 downto 54);
    -- logger for split-operator slice_1404_inst flow-through 
    process(addr2_1405) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:slice_1404_inst:flowthrough inputs: " & " cmd_1_1389 = "& Convert_SLV_To_Hex_String(cmd_1_1389) & " outputs:" & " addr2_1405= "  & Convert_SLV_To_Hex_String(addr2_1405));
      --
    end process; 
    -- flow-through slice operator slice_1404_inst
    addr2_1405 <= cmd_1_1389(53 downto 46);
    -- logger for split-operator slice_1408_inst flow-through 
    process(valid_w_1409) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:slice_1408_inst:flowthrough inputs: " & " cmd_1_1389 = "& Convert_SLV_To_Hex_String(cmd_1_1389) & " outputs:" & " valid_w_1409= "  & Convert_SLV_To_Hex_String(valid_w_1409));
      --
    end process; 
    -- flow-through slice operator slice_1408_inst
    valid_w_1409 <= cmd_1_1389(40 downto 40);
    -- logger for split-operator slice_1412_inst flow-through 
    process(addr_w_1413) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:slice_1412_inst:flowthrough inputs: " & " cmd_1_1389 = "& Convert_SLV_To_Hex_String(cmd_1_1389) & " outputs:" & " addr_w_1413= "  & Convert_SLV_To_Hex_String(addr_w_1413));
      --
    end process; 
    -- flow-through slice operator slice_1412_inst
    addr_w_1413 <= cmd_1_1389(39 downto 32);
    -- logger for split-operator slice_1416_inst flow-through 
    process(data_to_be_written_1417) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:slice_1416_inst:flowthrough inputs: " & " cmd_1_1389 = "& Convert_SLV_To_Hex_String(cmd_1_1389) & " outputs:" & " data_to_be_written_1417= "  & Convert_SLV_To_Hex_String(data_to_be_written_1417));
      --
    end process; 
    -- flow-through slice operator slice_1416_inst
    data_to_be_written_1417 <= cmd_1_1389(31 downto 0);
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1385_branch_req_0," req0 do_while_stmt_1385_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1385_branch_ack_0," ack0 do_while_stmt_1385_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1385_branch_ack_1," ack1 do_while_stmt_1385_branch");
    do_while_stmt_1385_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1435_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1385_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1385_branch_req_0,
          ack0 => do_while_stmt_1385_branch_ack_0,
          ack1 => do_while_stmt_1385_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_accessReg_request_1388_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_accessReg_request_1388_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:RPIPE_accessReg_request_1388_inst:started:   PipeRead from accessReg_request inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_accessReg_request_1388_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:RPIPE_accessReg_request_1388_inst:finished:  outputs: " & " cmd_1_1389= "  & Convert_SLV_To_Hex_String(cmd_1_1389));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_accessReg_request_1388_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_accessReg_request_1388_inst_req_0;
      RPIPE_accessReg_request_1388_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_accessReg_request_1388_inst_req_1;
      RPIPE_accessReg_request_1388_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      cmd_1_1389 <= data_out(63 downto 0);
      accessReg_request_read_0_gI: SplitGuardInterface generic map(name => "accessReg_request_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      accessReg_request_read_0: InputPortRevised -- 
        generic map ( name => "accessReg_request_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => accessReg_request_pipe_read_req(0),
          oack => accessReg_request_pipe_read_ack(0),
          odata => accessReg_request_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_accessReg_response1_1428_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_accessReg_response1_1428_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:WPIPE_accessReg_response1_1428_inst:started:   PipeWrite to accessReg_response1 inputs: " & " rdata1_1427 = "& Convert_SLV_To_Hex_String(rdata1_1427));
          --
        end if; 
        if WPIPE_accessReg_response1_1428_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:WPIPE_accessReg_response1_1428_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_accessReg_response1_1428_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_accessReg_response1_1428_inst_req_0;
      WPIPE_accessReg_response1_1428_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_accessReg_response1_1428_inst_req_1;
      WPIPE_accessReg_response1_1428_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= rdata1_1427;
      accessReg_response1_write_0_gI: SplitGuardInterface generic map(name => "accessReg_response1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      accessReg_response1_write_0: OutputPortRevised -- 
        generic map ( name => "accessReg_response1", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => accessReg_response1_pipe_write_req(0),
          oack => accessReg_response1_pipe_write_ack(0),
          odata => accessReg_response1_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_accessReg_response2_1431_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_accessReg_response2_1431_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:WPIPE_accessReg_response2_1431_inst:started:   PipeWrite to accessReg_response2 inputs: " & " rdata2_1427 = "& Convert_SLV_To_Hex_String(rdata2_1427));
          --
        end if; 
        if WPIPE_accessReg_response2_1431_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:WPIPE_accessReg_response2_1431_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_accessReg_response2_1431_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_accessReg_response2_1431_inst_req_0;
      WPIPE_accessReg_response2_1431_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_accessReg_response2_1431_inst_req_1;
      WPIPE_accessReg_response2_1431_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= rdata2_1427;
      accessReg_response2_write_1_gI: SplitGuardInterface generic map(name => "accessReg_response2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      accessReg_response2_write_1: OutputPortRevised -- 
        generic map ( name => "accessReg_response2", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => accessReg_response2_pipe_write_req(0),
          oack => accessReg_response2_pipe_write_ack(0),
          odata => accessReg_response2_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator call_stmt_1427_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1427_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:call_stmt_1427_call:started:  Call to module accessReg inputs: " & " valid_1_1393 = "& Convert_SLV_To_Hex_String(valid_1_1393) & " addr1_1397 = "& Convert_SLV_To_Hex_String(addr1_1397) & " valid_2_1401 = "& Convert_SLV_To_Hex_String(valid_2_1401) & " addr2_1405 = "& Convert_SLV_To_Hex_String(addr2_1405) & " valid_w_1409 = "& Convert_SLV_To_Hex_String(valid_w_1409) & " addr_w_1413 = "& Convert_SLV_To_Hex_String(addr_w_1413) & " data_to_be_written_1417 = "& Convert_SLV_To_Hex_String(data_to_be_written_1417));
          --
        end if; 
        if call_stmt_1427_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:regAccessDaemon:DP:call_stmt_1427_call:finished:  outputs: " & " rdata1_1427= "  & Convert_SLV_To_Hex_String(rdata1_1427) & " rdata2_1427= "  & Convert_SLV_To_Hex_String(rdata2_1427));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1427_call 
    accessReg_call_group_0: Block -- 
      signal data_in: std_logic_vector(58 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 7);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1427_call_req_0;
      call_stmt_1427_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1427_call_req_1;
      call_stmt_1427_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessReg_call_group_0_gI: SplitGuardInterface generic map(name => "accessReg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= valid_1_1393 & addr1_1397 & valid_2_1401 & addr2_1405 & valid_w_1409 & addr_w_1413 & data_to_be_written_1417;
      rdata1_1427 <= data_out(63 downto 32);
      rdata2_1427 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 59,
        owidth => 59,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessReg_call_reqs(0),
          ackR => accessReg_call_acks(0),
          dataR => accessReg_call_data(58 downto 0),
          tagR => accessReg_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessReg_return_acks(0), -- cross-over
          ackL => accessReg_return_reqs(0), -- cross-over
          dataL => accessReg_return_data(63 downto 0),
          tagL => accessReg_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end regAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity scoreBoard_Volatile is -- 
  port ( -- 
    clk, reset: in std_logic; 
    ifetch_state : in  std_logic_vector(9 downto 0);
    icache_state : in  std_logic_vector(9 downto 0);
    idecode_state : in  std_logic_vector(41 downto 0);
    iregfile_state : in  std_logic_vector(41 downto 0);
    iexec_state : in  std_logic_vector(105 downto 0);
    dcache_state : in  std_logic_vector(138 downto 0);
    iretire_state : in  std_logic_vector(138 downto 0);
    ifetch_actions : out  std_logic_vector(9 downto 0);
    icache_actions : out  std_logic_vector(9 downto 0);
    idecode_actions : out  std_logic_vector(41 downto 0);
    iregfile_actions : out  std_logic_vector(4 downto 0);
    iexec_actions : out  std_logic_vector(3 downto 0);
    dcache_actions : out  std_logic_vector(2 downto 0);
    ex_Unconditional_JUMP : out  std_logic_vector(0 downto 0);
    is_Branch_Hazard : out  std_logic_vector(0 downto 0);
    flush_ifetch : out  std_logic_vector(0 downto 0);
    flush_icache : out  std_logic_vector(0 downto 0);
    flush_idecode : out  std_logic_vector(0 downto 0);
    flush_reg : out  std_logic_vector(0 downto 0);
    flush_iexec : out  std_logic_vector(0 downto 0);
    flush_dcache : out  std_logic_vector(0 downto 0);
    stall_first_4 : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity scoreBoard_Volatile;
architecture scoreBoard_Volatile_arch of scoreBoard_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(488-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal ifetch_state_buffer :  std_logic_vector(9 downto 0);
  signal icache_state_buffer :  std_logic_vector(9 downto 0);
  signal idecode_state_buffer :  std_logic_vector(41 downto 0);
  signal iregfile_state_buffer :  std_logic_vector(41 downto 0);
  signal iexec_state_buffer :  std_logic_vector(105 downto 0);
  signal dcache_state_buffer :  std_logic_vector(138 downto 0);
  signal iretire_state_buffer :  std_logic_vector(138 downto 0);
  -- output port buffer signals
  signal ifetch_actions_buffer :  std_logic_vector(9 downto 0);
  signal icache_actions_buffer :  std_logic_vector(9 downto 0);
  signal idecode_actions_buffer :  std_logic_vector(41 downto 0);
  signal iregfile_actions_buffer :  std_logic_vector(4 downto 0);
  signal iexec_actions_buffer :  std_logic_vector(3 downto 0);
  signal dcache_actions_buffer :  std_logic_vector(2 downto 0);
  signal ex_Unconditional_JUMP_buffer :  std_logic_vector(0 downto 0);
  signal is_Branch_Hazard_buffer :  std_logic_vector(0 downto 0);
  signal flush_ifetch_buffer :  std_logic_vector(0 downto 0);
  signal flush_icache_buffer :  std_logic_vector(0 downto 0);
  signal flush_idecode_buffer :  std_logic_vector(0 downto 0);
  signal flush_reg_buffer :  std_logic_vector(0 downto 0);
  signal flush_iexec_buffer :  std_logic_vector(0 downto 0);
  signal flush_dcache_buffer :  std_logic_vector(0 downto 0);
  signal stall_first_4_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  ifetch_state_buffer <= ifetch_state;
  icache_state_buffer <= icache_state;
  idecode_state_buffer <= idecode_state;
  iregfile_state_buffer <= iregfile_state;
  iexec_state_buffer <= iexec_state;
  dcache_state_buffer <= dcache_state;
  iretire_state_buffer <= iretire_state;
  -- output handling  -------------------------------------------------------
  ifetch_actions <= ifetch_actions_buffer;
  icache_actions <= icache_actions_buffer;
  idecode_actions <= idecode_actions_buffer;
  iregfile_actions <= iregfile_actions_buffer;
  iexec_actions <= iexec_actions_buffer;
  dcache_actions <= dcache_actions_buffer;
  ex_Unconditional_JUMP <= ex_Unconditional_JUMP_buffer;
  is_Branch_Hazard <= is_Branch_Hazard_buffer;
  flush_ifetch <= flush_ifetch_buffer;
  flush_icache <= flush_icache_buffer;
  flush_idecode <= flush_idecode_buffer;
  flush_reg <= flush_reg_buffer;
  flush_iexec <= flush_iexec_buffer;
  flush_dcache <= flush_dcache_buffer;
  stall_first_4 <= stall_first_4_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_785_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_797_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u1_u2_887_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_892_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_898_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_901_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_915_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u3_889_wire : std_logic_vector(2 downto 0);
    signal EQ_u1_u1_635_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_644_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_714_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_723_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_732_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_741_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_762_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_771_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_803_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_806_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_812_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_815_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_821_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_824_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_830_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_833_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_839_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_842_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_846_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_558_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_561_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_586_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_589_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_593_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_597_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_600_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_604_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_609_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_612_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_616_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_620_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_623_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_627_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_638_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_647_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_665_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_668_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_672_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_676_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_679_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_683_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_688_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_691_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_695_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_699_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_702_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_706_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_717_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_726_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_735_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_744_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_765_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_774_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_780_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_783_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_788_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_792_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_795_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_868_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_876_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_907_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_784_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_789_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_590_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_594_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_601_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_605_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_606_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_613_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_617_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_624_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_628_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_629_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_669_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_673_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_680_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_684_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_685_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_692_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_696_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_703_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_707_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_708_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_796_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_843_wire : std_logic_vector(0 downto 0);
    signal R_ADD_603_wire_constant : std_logic_vector(7 downto 0);
    signal R_ADD_682_wire_constant : std_logic_vector(7 downto 0);
    signal R_CALL_557_wire_constant : std_logic_vector(7 downto 0);
    signal R_CALL_622_wire_constant : std_logic_vector(7 downto 0);
    signal R_CALL_701_wire_constant : std_logic_vector(7 downto 0);
    signal R_CMP_626_wire_constant : std_logic_vector(7 downto 0);
    signal R_CMP_705_wire_constant : std_logic_vector(7 downto 0);
    signal R_JMP_560_wire_constant : std_logic_vector(7 downto 0);
    signal R_LOAD_588_wire_constant : std_logic_vector(7 downto 0);
    signal R_LOAD_667_wire_constant : std_logic_vector(7 downto 0);
    signal R_LOAD_779_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_AND_592_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_AND_671_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_OR_596_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_OR_675_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SLL_611_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SLL_690_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SRA_619_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SRA_698_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SRL_615_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_SRL_694_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_XNOR_599_wire_constant : std_logic_vector(7 downto 0);
    signal R_L_XNOR_678_wire_constant : std_logic_vector(7 downto 0);
    signal R_SBIR_585_wire_constant : std_logic_vector(7 downto 0);
    signal R_SBIR_664_wire_constant : std_logic_vector(7 downto 0);
    signal R_STORE_787_wire_constant : std_logic_vector(7 downto 0);
    signal R_STORE_906_wire_constant : std_logic_vector(7 downto 0);
    signal R_SUB_608_wire_constant : std_logic_vector(7 downto 0);
    signal R_SUB_687_wire_constant : std_logic_vector(7 downto 0);
    signal R_one_1_634_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_643_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_713_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_722_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_731_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_740_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_761_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_770_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_802_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_805_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_811_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_814_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_820_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_823_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_829_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_832_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_838_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_841_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_845_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_870_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_878_wire_constant : std_logic_vector(0 downto 0);
    signal R_one_1_909_wire_constant : std_logic_vector(0 downto 0);
    signal R_zero_1_869_wire_constant : std_logic_vector(0 downto 0);
    signal R_zero_1_877_wire_constant : std_logic_vector(0 downto 0);
    signal R_zero_1_908_wire_constant : std_logic_vector(0 downto 0);
    signal R_zero_8_782_wire_constant : std_logic_vector(7 downto 0);
    signal dcache_opcode_570 : std_logic_vector(7 downto 0);
    signal dcache_rd_582 : std_logic_vector(7 downto 0);
    signal dcache_rs1_imm_574 : std_logic_vector(7 downto 0);
    signal dcache_rs2_578 : std_logic_vector(7 downto 0);
    signal dcache_state_reg_write_631 : std_logic_vector(0 downto 0);
    signal dcache_to_ex_rs1_imm_640 : std_logic_vector(0 downto 0);
    signal dcache_to_ex_rs2_649 : std_logic_vector(0 downto 0);
    signal ex_opcode_542 : std_logic_vector(7 downto 0);
    signal ex_rd_554 : std_logic_vector(7 downto 0);
    signal ex_rs1_imm_546 : std_logic_vector(7 downto 0);
    signal ex_rs2_550 : std_logic_vector(7 downto 0);
    signal iregfile_opcode_750 : std_logic_vector(7 downto 0);
    signal iregfile_rs1_imm_754 : std_logic_vector(7 downto 0);
    signal iregfile_rs2_758 : std_logic_vector(7 downto 0);
    signal iregfile_state_opcode_864 : std_logic_vector(7 downto 0);
    signal iretire_opcode_653 : std_logic_vector(7 downto 0);
    signal iretire_rd_661 : std_logic_vector(7 downto 0);
    signal iretire_rs1_imm_657 : std_logic_vector(7 downto 0);
    signal iretire_state_reg_write_710 : std_logic_vector(0 downto 0);
    signal iretire_state_to_dcache_addr_737 : std_logic_vector(0 downto 0);
    signal iretire_state_to_dcache_memData_746 : std_logic_vector(0 downto 0);
    signal iretire_state_to_ex_rs1_imm_719 : std_logic_vector(0 downto 0);
    signal iretire_state_to_ex_rs2_728 : std_logic_vector(0 downto 0);
    signal iretire_state_to_rs1_imm_767 : std_logic_vector(0 downto 0);
    signal iretire_state_to_rs2_776 : std_logic_vector(0 downto 0);
    signal is_Branch_538 : std_logic_vector(0 downto 0);
    signal konst_867_wire_constant : std_logic_vector(7 downto 0);
    signal konst_875_wire_constant : std_logic_vector(7 downto 0);
    signal memWrite_911 : std_logic_vector(0 downto 0);
    signal reg_valid_read1_872 : std_logic_vector(0 downto 0);
    signal reg_valid_read2_880 : std_logic_vector(0 downto 0);
    signal reg_valid_write_883 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ADD_603_wire_constant <= "00001001";
    R_ADD_682_wire_constant <= "00001001";
    R_CALL_557_wire_constant <= "00010000";
    R_CALL_622_wire_constant <= "00010000";
    R_CALL_701_wire_constant <= "00010000";
    R_CMP_626_wire_constant <= "00010010";
    R_CMP_705_wire_constant <= "00010010";
    R_JMP_560_wire_constant <= "00010001";
    R_LOAD_588_wire_constant <= "00000011";
    R_LOAD_667_wire_constant <= "00000011";
    R_LOAD_779_wire_constant <= "00000011";
    R_L_AND_592_wire_constant <= "00000101";
    R_L_AND_671_wire_constant <= "00000101";
    R_L_OR_596_wire_constant <= "00000110";
    R_L_OR_675_wire_constant <= "00000110";
    R_L_SLL_611_wire_constant <= "00001011";
    R_L_SLL_690_wire_constant <= "00001011";
    R_L_SRA_619_wire_constant <= "00001101";
    R_L_SRA_698_wire_constant <= "00001101";
    R_L_SRL_615_wire_constant <= "00001100";
    R_L_SRL_694_wire_constant <= "00001100";
    R_L_XNOR_599_wire_constant <= "00000111";
    R_L_XNOR_678_wire_constant <= "00000111";
    R_SBIR_585_wire_constant <= "00000010";
    R_SBIR_664_wire_constant <= "00000010";
    R_STORE_787_wire_constant <= "00000100";
    R_STORE_906_wire_constant <= "00000100";
    R_SUB_608_wire_constant <= "00001010";
    R_SUB_687_wire_constant <= "00001010";
    R_one_1_634_wire_constant <= "1";
    R_one_1_643_wire_constant <= "1";
    R_one_1_713_wire_constant <= "1";
    R_one_1_722_wire_constant <= "1";
    R_one_1_731_wire_constant <= "1";
    R_one_1_740_wire_constant <= "1";
    R_one_1_761_wire_constant <= "1";
    R_one_1_770_wire_constant <= "1";
    R_one_1_802_wire_constant <= "1";
    R_one_1_805_wire_constant <= "1";
    R_one_1_811_wire_constant <= "1";
    R_one_1_814_wire_constant <= "1";
    R_one_1_820_wire_constant <= "1";
    R_one_1_823_wire_constant <= "1";
    R_one_1_829_wire_constant <= "1";
    R_one_1_832_wire_constant <= "1";
    R_one_1_838_wire_constant <= "1";
    R_one_1_841_wire_constant <= "1";
    R_one_1_845_wire_constant <= "1";
    R_one_1_870_wire_constant <= "1";
    R_one_1_878_wire_constant <= "1";
    R_one_1_909_wire_constant <= "1";
    R_zero_1_869_wire_constant <= "0";
    R_zero_1_877_wire_constant <= "0";
    R_zero_1_908_wire_constant <= "0";
    R_zero_8_782_wire_constant <= "00000000";
    konst_867_wire_constant <= "00000000";
    konst_875_wire_constant <= "00000000";
    -- logger for split-operator MUX_871_inst flow-through 
    process(reg_valid_read1_872) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:MUX_871_inst:flowthrough inputs: " & " EQ_u8_u1_868_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_868_wire) & " R_zero_1_869_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_1_869_wire_constant) & " R_one_1_870_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_870_wire_constant) & " outputs:" & " reg_valid_read1_872= "  & Convert_SLV_To_Hex_String(reg_valid_read1_872));
      --
    end process; 
    -- flow-through select operator MUX_871_inst
    reg_valid_read1_872 <= R_zero_1_869_wire_constant when (EQ_u8_u1_868_wire(0) /=  '0') else R_one_1_870_wire_constant;
    -- logger for split-operator MUX_879_inst flow-through 
    process(reg_valid_read2_880) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:MUX_879_inst:flowthrough inputs: " & " EQ_u8_u1_876_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_876_wire) & " R_zero_1_877_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_1_877_wire_constant) & " R_one_1_878_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_878_wire_constant) & " outputs:" & " reg_valid_read2_880= "  & Convert_SLV_To_Hex_String(reg_valid_read2_880));
      --
    end process; 
    -- flow-through select operator MUX_879_inst
    reg_valid_read2_880 <= R_zero_1_877_wire_constant when (EQ_u8_u1_876_wire(0) /=  '0') else R_one_1_878_wire_constant;
    -- logger for split-operator MUX_910_inst flow-through 
    process(memWrite_911) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:MUX_910_inst:flowthrough inputs: " & " EQ_u8_u1_907_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_907_wire) & " R_zero_1_908_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_1_908_wire_constant) & " R_one_1_909_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_909_wire_constant) & " outputs:" & " memWrite_911= "  & Convert_SLV_To_Hex_String(memWrite_911));
      --
    end process; 
    -- flow-through select operator MUX_910_inst
    memWrite_911 <= R_zero_1_908_wire_constant when (EQ_u8_u1_907_wire(0) /=  '0') else R_one_1_909_wire_constant;
    -- logger for split-operator slice_537_inst flow-through 
    process(is_Branch_538) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_537_inst:flowthrough inputs: " & " dcache_state_buffer = "& Convert_SLV_To_Hex_String(dcache_state_buffer) & " outputs:" & " is_Branch_538= "  & Convert_SLV_To_Hex_String(is_Branch_538));
      --
    end process; 
    -- flow-through slice operator slice_537_inst
    is_Branch_538 <= dcache_state_buffer(10 downto 10);
    -- logger for split-operator slice_541_inst flow-through 
    process(ex_opcode_542) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_541_inst:flowthrough inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer) & " outputs:" & " ex_opcode_542= "  & Convert_SLV_To_Hex_String(ex_opcode_542));
      --
    end process; 
    -- flow-through slice operator slice_541_inst
    ex_opcode_542 <= iexec_state_buffer(105 downto 98);
    -- logger for split-operator slice_545_inst flow-through 
    process(ex_rs1_imm_546) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_545_inst:flowthrough inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer) & " outputs:" & " ex_rs1_imm_546= "  & Convert_SLV_To_Hex_String(ex_rs1_imm_546));
      --
    end process; 
    -- flow-through slice operator slice_545_inst
    ex_rs1_imm_546 <= iexec_state_buffer(97 downto 90);
    -- logger for split-operator slice_549_inst flow-through 
    process(ex_rs2_550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_549_inst:flowthrough inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer) & " outputs:" & " ex_rs2_550= "  & Convert_SLV_To_Hex_String(ex_rs2_550));
      --
    end process; 
    -- flow-through slice operator slice_549_inst
    ex_rs2_550 <= iexec_state_buffer(89 downto 82);
    -- logger for split-operator slice_553_inst flow-through 
    process(ex_rd_554) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_553_inst:flowthrough inputs: " & " iexec_state_buffer = "& Convert_SLV_To_Hex_String(iexec_state_buffer) & " outputs:" & " ex_rd_554= "  & Convert_SLV_To_Hex_String(ex_rd_554));
      --
    end process; 
    -- flow-through slice operator slice_553_inst
    ex_rd_554 <= iexec_state_buffer(81 downto 74);
    -- logger for split-operator slice_569_inst flow-through 
    process(dcache_opcode_570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_569_inst:flowthrough inputs: " & " dcache_state_buffer = "& Convert_SLV_To_Hex_String(dcache_state_buffer) & " outputs:" & " dcache_opcode_570= "  & Convert_SLV_To_Hex_String(dcache_opcode_570));
      --
    end process; 
    -- flow-through slice operator slice_569_inst
    dcache_opcode_570 <= dcache_state_buffer(138 downto 131);
    -- logger for split-operator slice_573_inst flow-through 
    process(dcache_rs1_imm_574) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_573_inst:flowthrough inputs: " & " dcache_state_buffer = "& Convert_SLV_To_Hex_String(dcache_state_buffer) & " outputs:" & " dcache_rs1_imm_574= "  & Convert_SLV_To_Hex_String(dcache_rs1_imm_574));
      --
    end process; 
    -- flow-through slice operator slice_573_inst
    dcache_rs1_imm_574 <= dcache_state_buffer(130 downto 123);
    -- logger for split-operator slice_577_inst flow-through 
    process(dcache_rs2_578) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_577_inst:flowthrough inputs: " & " dcache_state_buffer = "& Convert_SLV_To_Hex_String(dcache_state_buffer) & " outputs:" & " dcache_rs2_578= "  & Convert_SLV_To_Hex_String(dcache_rs2_578));
      --
    end process; 
    -- flow-through slice operator slice_577_inst
    dcache_rs2_578 <= dcache_state_buffer(122 downto 115);
    -- logger for split-operator slice_581_inst flow-through 
    process(dcache_rd_582) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_581_inst:flowthrough inputs: " & " dcache_state_buffer = "& Convert_SLV_To_Hex_String(dcache_state_buffer) & " outputs:" & " dcache_rd_582= "  & Convert_SLV_To_Hex_String(dcache_rd_582));
      --
    end process; 
    -- flow-through slice operator slice_581_inst
    dcache_rd_582 <= dcache_state_buffer(114 downto 107);
    -- logger for split-operator slice_652_inst flow-through 
    process(iretire_opcode_653) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_652_inst:flowthrough inputs: " & " iretire_state_buffer = "& Convert_SLV_To_Hex_String(iretire_state_buffer) & " outputs:" & " iretire_opcode_653= "  & Convert_SLV_To_Hex_String(iretire_opcode_653));
      --
    end process; 
    -- flow-through slice operator slice_652_inst
    iretire_opcode_653 <= iretire_state_buffer(138 downto 131);
    -- logger for split-operator slice_656_inst flow-through 
    process(iretire_rs1_imm_657) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_656_inst:flowthrough inputs: " & " iretire_state_buffer = "& Convert_SLV_To_Hex_String(iretire_state_buffer) & " outputs:" & " iretire_rs1_imm_657= "  & Convert_SLV_To_Hex_String(iretire_rs1_imm_657));
      --
    end process; 
    -- flow-through slice operator slice_656_inst
    iretire_rs1_imm_657 <= iretire_state_buffer(130 downto 123);
    -- logger for split-operator slice_660_inst flow-through 
    process(iretire_rd_661) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_660_inst:flowthrough inputs: " & " iretire_state_buffer = "& Convert_SLV_To_Hex_String(iretire_state_buffer) & " outputs:" & " iretire_rd_661= "  & Convert_SLV_To_Hex_String(iretire_rd_661));
      --
    end process; 
    -- flow-through slice operator slice_660_inst
    iretire_rd_661 <= iretire_state_buffer(114 downto 107);
    -- logger for split-operator slice_749_inst flow-through 
    process(iregfile_opcode_750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_749_inst:flowthrough inputs: " & " iregfile_state_buffer = "& Convert_SLV_To_Hex_String(iregfile_state_buffer) & " outputs:" & " iregfile_opcode_750= "  & Convert_SLV_To_Hex_String(iregfile_opcode_750));
      --
    end process; 
    -- flow-through slice operator slice_749_inst
    iregfile_opcode_750 <= iregfile_state_buffer(41 downto 34);
    -- logger for split-operator slice_753_inst flow-through 
    process(iregfile_rs1_imm_754) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_753_inst:flowthrough inputs: " & " iregfile_state_buffer = "& Convert_SLV_To_Hex_String(iregfile_state_buffer) & " outputs:" & " iregfile_rs1_imm_754= "  & Convert_SLV_To_Hex_String(iregfile_rs1_imm_754));
      --
    end process; 
    -- flow-through slice operator slice_753_inst
    iregfile_rs1_imm_754 <= iregfile_state_buffer(33 downto 26);
    -- logger for split-operator slice_757_inst flow-through 
    process(iregfile_rs2_758) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_757_inst:flowthrough inputs: " & " iregfile_state_buffer = "& Convert_SLV_To_Hex_String(iregfile_state_buffer) & " outputs:" & " iregfile_rs2_758= "  & Convert_SLV_To_Hex_String(iregfile_rs2_758));
      --
    end process; 
    -- flow-through slice operator slice_757_inst
    iregfile_rs2_758 <= iregfile_state_buffer(25 downto 18);
    -- logger for split-operator slice_863_inst flow-through 
    process(iregfile_state_opcode_864) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:slice_863_inst:flowthrough inputs: " & " iregfile_state_buffer = "& Convert_SLV_To_Hex_String(iregfile_state_buffer) & " outputs:" & " iregfile_state_opcode_864= "  & Convert_SLV_To_Hex_String(iregfile_state_opcode_864));
      --
    end process; 
    -- flow-through slice operator slice_863_inst
    iregfile_state_opcode_864 <= iregfile_state_buffer(41 downto 34);
    -- logger for split-operator W_flush_dcache_849_inst flow-through 
    process(flush_dcache_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:W_flush_dcache_849_inst:flowthrough inputs: " & " is_Branch_538 = "& Convert_SLV_To_Hex_String(is_Branch_538) & " outputs:" & " flush_dcache_buffer= "  & Convert_SLV_To_Hex_String(flush_dcache_buffer));
      --
    end process; 
    -- interlock W_flush_dcache_849_inst
    process(is_Branch_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := is_Branch_538(0 downto 0);
      flush_dcache_buffer <= tmp_var; -- 
    end process;
    -- logger for split-operator W_icache_actions_855_inst flow-through 
    process(icache_actions_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:W_icache_actions_855_inst:flowthrough inputs: " & " icache_state_buffer = "& Convert_SLV_To_Hex_String(icache_state_buffer) & " outputs:" & " icache_actions_buffer= "  & Convert_SLV_To_Hex_String(icache_actions_buffer));
      --
    end process; 
    -- interlock W_icache_actions_855_inst
    process(icache_state_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 9 downto 0) := icache_state_buffer(9 downto 0);
      icache_actions_buffer <= tmp_var; -- 
    end process;
    -- logger for split-operator W_idecode_actions_858_inst flow-through 
    process(idecode_actions_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:W_idecode_actions_858_inst:flowthrough inputs: " & " idecode_state_buffer = "& Convert_SLV_To_Hex_String(idecode_state_buffer) & " outputs:" & " idecode_actions_buffer= "  & Convert_SLV_To_Hex_String(idecode_actions_buffer));
      --
    end process; 
    -- interlock W_idecode_actions_858_inst
    process(idecode_state_buffer) -- 
      variable tmp_var : std_logic_vector(41 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 41 downto 0) := idecode_state_buffer(41 downto 0);
      idecode_actions_buffer <= tmp_var; -- 
    end process;
    -- logger for split-operator W_ifetch_actions_852_inst flow-through 
    process(ifetch_actions_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:W_ifetch_actions_852_inst:flowthrough inputs: " & " ifetch_state_buffer = "& Convert_SLV_To_Hex_String(ifetch_state_buffer) & " outputs:" & " ifetch_actions_buffer= "  & Convert_SLV_To_Hex_String(ifetch_actions_buffer));
      --
    end process; 
    -- interlock W_ifetch_actions_852_inst
    process(ifetch_state_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 9 downto 0) := ifetch_state_buffer(9 downto 0);
      ifetch_actions_buffer <= tmp_var; -- 
    end process;
    -- logger for split-operator W_is_Branch_Hazard_564_inst flow-through 
    process(is_Branch_Hazard_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:W_is_Branch_Hazard_564_inst:flowthrough inputs: " & " is_Branch_538 = "& Convert_SLV_To_Hex_String(is_Branch_538) & " outputs:" & " is_Branch_Hazard_buffer= "  & Convert_SLV_To_Hex_String(is_Branch_Hazard_buffer));
      --
    end process; 
    -- interlock W_is_Branch_Hazard_564_inst
    process(is_Branch_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := is_Branch_538(0 downto 0);
      is_Branch_Hazard_buffer <= tmp_var; -- 
    end process;
    -- logger for split-operator W_reg_valid_write_881_inst flow-through 
    process(reg_valid_write_883) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:W_reg_valid_write_881_inst:flowthrough inputs: " & " iretire_state_reg_write_710 = "& Convert_SLV_To_Hex_String(iretire_state_reg_write_710) & " outputs:" & " reg_valid_write_883= "  & Convert_SLV_To_Hex_String(reg_valid_write_883));
      --
    end process; 
    -- interlock W_reg_valid_write_881_inst
    process(iretire_state_reg_write_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := iretire_state_reg_write_710(0 downto 0);
      reg_valid_write_883 <= tmp_var; -- 
    end process;
    -- logger for split-operator AND_u1_u1_639_inst flow-through 
    process(dcache_to_ex_rs1_imm_640) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_639_inst:flowthrough inputs: " & " EQ_u1_u1_635_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_635_wire) & " EQ_u8_u1_638_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_638_wire) & " outputs:" & " dcache_to_ex_rs1_imm_640= "  & Convert_SLV_To_Hex_String(dcache_to_ex_rs1_imm_640));
      --
    end process; 
    -- binary operator AND_u1_u1_639_inst
    process(EQ_u1_u1_635_wire, EQ_u8_u1_638_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_635_wire, EQ_u8_u1_638_wire, tmp_var);
      dcache_to_ex_rs1_imm_640 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_648_inst flow-through 
    process(dcache_to_ex_rs2_649) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_648_inst:flowthrough inputs: " & " EQ_u1_u1_644_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_644_wire) & " EQ_u8_u1_647_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_647_wire) & " outputs:" & " dcache_to_ex_rs2_649= "  & Convert_SLV_To_Hex_String(dcache_to_ex_rs2_649));
      --
    end process; 
    -- binary operator AND_u1_u1_648_inst
    process(EQ_u1_u1_644_wire, EQ_u8_u1_647_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_644_wire, EQ_u8_u1_647_wire, tmp_var);
      dcache_to_ex_rs2_649 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_718_inst flow-through 
    process(iretire_state_to_ex_rs1_imm_719) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_718_inst:flowthrough inputs: " & " EQ_u1_u1_714_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_714_wire) & " EQ_u8_u1_717_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_717_wire) & " outputs:" & " iretire_state_to_ex_rs1_imm_719= "  & Convert_SLV_To_Hex_String(iretire_state_to_ex_rs1_imm_719));
      --
    end process; 
    -- binary operator AND_u1_u1_718_inst
    process(EQ_u1_u1_714_wire, EQ_u8_u1_717_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_714_wire, EQ_u8_u1_717_wire, tmp_var);
      iretire_state_to_ex_rs1_imm_719 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_727_inst flow-through 
    process(iretire_state_to_ex_rs2_728) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_727_inst:flowthrough inputs: " & " EQ_u1_u1_723_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_723_wire) & " EQ_u8_u1_726_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_726_wire) & " outputs:" & " iretire_state_to_ex_rs2_728= "  & Convert_SLV_To_Hex_String(iretire_state_to_ex_rs2_728));
      --
    end process; 
    -- binary operator AND_u1_u1_727_inst
    process(EQ_u1_u1_723_wire, EQ_u8_u1_726_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_723_wire, EQ_u8_u1_726_wire, tmp_var);
      iretire_state_to_ex_rs2_728 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_736_inst flow-through 
    process(iretire_state_to_dcache_addr_737) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_736_inst:flowthrough inputs: " & " EQ_u1_u1_732_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_732_wire) & " EQ_u8_u1_735_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_735_wire) & " outputs:" & " iretire_state_to_dcache_addr_737= "  & Convert_SLV_To_Hex_String(iretire_state_to_dcache_addr_737));
      --
    end process; 
    -- binary operator AND_u1_u1_736_inst
    process(EQ_u1_u1_732_wire, EQ_u8_u1_735_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_732_wire, EQ_u8_u1_735_wire, tmp_var);
      iretire_state_to_dcache_addr_737 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_745_inst flow-through 
    process(iretire_state_to_dcache_memData_746) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_745_inst:flowthrough inputs: " & " EQ_u1_u1_741_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_741_wire) & " EQ_u8_u1_744_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_744_wire) & " outputs:" & " iretire_state_to_dcache_memData_746= "  & Convert_SLV_To_Hex_String(iretire_state_to_dcache_memData_746));
      --
    end process; 
    -- binary operator AND_u1_u1_745_inst
    process(EQ_u1_u1_741_wire, EQ_u8_u1_744_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_741_wire, EQ_u8_u1_744_wire, tmp_var);
      iretire_state_to_dcache_memData_746 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_766_inst flow-through 
    process(iretire_state_to_rs1_imm_767) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_766_inst:flowthrough inputs: " & " EQ_u1_u1_762_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_762_wire) & " EQ_u8_u1_765_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_765_wire) & " outputs:" & " iretire_state_to_rs1_imm_767= "  & Convert_SLV_To_Hex_String(iretire_state_to_rs1_imm_767));
      --
    end process; 
    -- binary operator AND_u1_u1_766_inst
    process(EQ_u1_u1_762_wire, EQ_u8_u1_765_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_762_wire, EQ_u8_u1_765_wire, tmp_var);
      iretire_state_to_rs1_imm_767 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_775_inst flow-through 
    process(iretire_state_to_rs2_776) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_775_inst:flowthrough inputs: " & " EQ_u1_u1_771_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_771_wire) & " EQ_u8_u1_774_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_774_wire) & " outputs:" & " iretire_state_to_rs2_776= "  & Convert_SLV_To_Hex_String(iretire_state_to_rs2_776));
      --
    end process; 
    -- binary operator AND_u1_u1_775_inst
    process(EQ_u1_u1_771_wire, EQ_u8_u1_774_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_771_wire, EQ_u8_u1_774_wire, tmp_var);
      iretire_state_to_rs2_776 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_785_inst flow-through 
    process(AND_u1_u1_785_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_785_inst:flowthrough inputs: " & " EQ_u8_u1_780_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_780_wire) & " NOT_u1_u1_784_wire = "& Convert_SLV_To_Hex_String(NOT_u1_u1_784_wire) & " outputs:" & " AND_u1_u1_785_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_785_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_785_inst
    process(EQ_u8_u1_780_wire, NOT_u1_u1_784_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u8_u1_780_wire, NOT_u1_u1_784_wire, tmp_var);
      AND_u1_u1_785_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_797_inst flow-through 
    process(AND_u1_u1_797_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_797_inst:flowthrough inputs: " & " NOT_u1_u1_789_wire = "& Convert_SLV_To_Hex_String(NOT_u1_u1_789_wire) & " OR_u1_u1_796_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_796_wire) & " outputs:" & " AND_u1_u1_797_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_797_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_797_inst
    process(NOT_u1_u1_789_wire, OR_u1_u1_796_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_789_wire, OR_u1_u1_796_wire, tmp_var);
      AND_u1_u1_797_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_798_inst flow-through 
    process(stall_first_4_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:AND_u1_u1_798_inst:flowthrough inputs: " & " AND_u1_u1_785_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_785_wire) & " AND_u1_u1_797_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_797_wire) & " outputs:" & " stall_first_4_buffer= "  & Convert_SLV_To_Hex_String(stall_first_4_buffer));
      --
    end process; 
    -- binary operator AND_u1_u1_798_inst
    process(AND_u1_u1_785_wire, AND_u1_u1_797_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_785_wire, AND_u1_u1_797_wire, tmp_var);
      stall_first_4_buffer <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u2_887_inst flow-through 
    process(CONCAT_u1_u2_887_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u1_u2_887_inst:flowthrough inputs: " & " reg_valid_read1_872 = "& Convert_SLV_To_Hex_String(reg_valid_read1_872) & " reg_valid_read2_880 = "& Convert_SLV_To_Hex_String(reg_valid_read2_880) & " outputs:" & " CONCAT_u1_u2_887_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u2_887_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u2_887_inst
    process(reg_valid_read1_872, reg_valid_read2_880) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(reg_valid_read1_872, reg_valid_read2_880, tmp_var);
      CONCAT_u1_u2_887_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u2_892_inst flow-through 
    process(CONCAT_u1_u2_892_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u1_u2_892_inst:flowthrough inputs: " & " iretire_state_to_rs1_imm_767 = "& Convert_SLV_To_Hex_String(iretire_state_to_rs1_imm_767) & " iretire_state_to_rs2_776 = "& Convert_SLV_To_Hex_String(iretire_state_to_rs2_776) & " outputs:" & " CONCAT_u1_u2_892_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u2_892_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u2_892_inst
    process(iretire_state_to_rs1_imm_767, iretire_state_to_rs2_776) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(iretire_state_to_rs1_imm_767, iretire_state_to_rs2_776, tmp_var);
      CONCAT_u1_u2_892_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u2_898_inst flow-through 
    process(CONCAT_u1_u2_898_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u1_u2_898_inst:flowthrough inputs: " & " dcache_to_ex_rs1_imm_640 = "& Convert_SLV_To_Hex_String(dcache_to_ex_rs1_imm_640) & " dcache_to_ex_rs2_649 = "& Convert_SLV_To_Hex_String(dcache_to_ex_rs2_649) & " outputs:" & " CONCAT_u1_u2_898_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u2_898_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u2_898_inst
    process(dcache_to_ex_rs1_imm_640, dcache_to_ex_rs2_649) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(dcache_to_ex_rs1_imm_640, dcache_to_ex_rs2_649, tmp_var);
      CONCAT_u1_u2_898_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u2_901_inst flow-through 
    process(CONCAT_u1_u2_901_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u1_u2_901_inst:flowthrough inputs: " & " iretire_state_to_ex_rs1_imm_719 = "& Convert_SLV_To_Hex_String(iretire_state_to_ex_rs1_imm_719) & " iretire_state_to_ex_rs2_728 = "& Convert_SLV_To_Hex_String(iretire_state_to_ex_rs2_728) & " outputs:" & " CONCAT_u1_u2_901_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u2_901_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u2_901_inst
    process(iretire_state_to_ex_rs1_imm_719, iretire_state_to_ex_rs2_728) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(iretire_state_to_ex_rs1_imm_719, iretire_state_to_ex_rs2_728, tmp_var);
      CONCAT_u1_u2_901_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u2_915_inst flow-through 
    process(CONCAT_u1_u2_915_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u1_u2_915_inst:flowthrough inputs: " & " memWrite_911 = "& Convert_SLV_To_Hex_String(memWrite_911) & " iretire_state_to_dcache_addr_737 = "& Convert_SLV_To_Hex_String(iretire_state_to_dcache_addr_737) & " outputs:" & " CONCAT_u1_u2_915_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u2_915_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u2_915_inst
    process(memWrite_911, iretire_state_to_dcache_addr_737) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(memWrite_911, iretire_state_to_dcache_addr_737, tmp_var);
      CONCAT_u1_u2_915_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u2_u3_889_inst flow-through 
    process(CONCAT_u2_u3_889_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u2_u3_889_inst:flowthrough inputs: " & " CONCAT_u1_u2_887_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u2_887_wire) & " reg_valid_write_883 = "& Convert_SLV_To_Hex_String(reg_valid_write_883) & " outputs:" & " CONCAT_u2_u3_889_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u2_u3_889_wire));
      --
    end process; 
    -- binary operator CONCAT_u2_u3_889_inst
    process(CONCAT_u1_u2_887_wire, reg_valid_write_883) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_887_wire, reg_valid_write_883, tmp_var);
      CONCAT_u2_u3_889_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u2_u3_917_inst flow-through 
    process(dcache_actions_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u2_u3_917_inst:flowthrough inputs: " & " CONCAT_u1_u2_915_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u2_915_wire) & " iretire_state_to_dcache_memData_746 = "& Convert_SLV_To_Hex_String(iretire_state_to_dcache_memData_746) & " outputs:" & " dcache_actions_buffer= "  & Convert_SLV_To_Hex_String(dcache_actions_buffer));
      --
    end process; 
    -- binary operator CONCAT_u2_u3_917_inst
    process(CONCAT_u1_u2_915_wire, iretire_state_to_dcache_memData_746) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_915_wire, iretire_state_to_dcache_memData_746, tmp_var);
      dcache_actions_buffer <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u2_u4_902_inst flow-through 
    process(iexec_actions_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u2_u4_902_inst:flowthrough inputs: " & " CONCAT_u1_u2_898_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u2_898_wire) & " CONCAT_u1_u2_901_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u2_901_wire) & " outputs:" & " iexec_actions_buffer= "  & Convert_SLV_To_Hex_String(iexec_actions_buffer));
      --
    end process; 
    -- binary operator CONCAT_u2_u4_902_inst
    process(CONCAT_u1_u2_898_wire, CONCAT_u1_u2_901_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_898_wire, CONCAT_u1_u2_901_wire, tmp_var);
      iexec_actions_buffer <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u3_u5_893_inst flow-through 
    process(iregfile_actions_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:CONCAT_u3_u5_893_inst:flowthrough inputs: " & " CONCAT_u2_u3_889_wire = "& Convert_SLV_To_Hex_String(CONCAT_u2_u3_889_wire) & " CONCAT_u1_u2_892_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u2_892_wire) & " outputs:" & " iregfile_actions_buffer= "  & Convert_SLV_To_Hex_String(iregfile_actions_buffer));
      --
    end process; 
    -- binary operator CONCAT_u3_u5_893_inst
    process(CONCAT_u2_u3_889_wire, CONCAT_u1_u2_892_wire) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u3_889_wire, CONCAT_u1_u2_892_wire, tmp_var);
      iregfile_actions_buffer <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_635_inst flow-through 
    process(EQ_u1_u1_635_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_635_inst:flowthrough inputs: " & " dcache_state_reg_write_631 = "& Convert_SLV_To_Hex_String(dcache_state_reg_write_631) & " R_one_1_634_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_634_wire_constant) & " outputs:" & " EQ_u1_u1_635_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_635_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_635_inst
    process(dcache_state_reg_write_631) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_state_reg_write_631, R_one_1_634_wire_constant, tmp_var);
      EQ_u1_u1_635_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_644_inst flow-through 
    process(EQ_u1_u1_644_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_644_inst:flowthrough inputs: " & " dcache_state_reg_write_631 = "& Convert_SLV_To_Hex_String(dcache_state_reg_write_631) & " R_one_1_643_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_643_wire_constant) & " outputs:" & " EQ_u1_u1_644_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_644_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_644_inst
    process(dcache_state_reg_write_631) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_state_reg_write_631, R_one_1_643_wire_constant, tmp_var);
      EQ_u1_u1_644_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_714_inst flow-through 
    process(EQ_u1_u1_714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_714_inst:flowthrough inputs: " & " iretire_state_reg_write_710 = "& Convert_SLV_To_Hex_String(iretire_state_reg_write_710) & " R_one_1_713_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_713_wire_constant) & " outputs:" & " EQ_u1_u1_714_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_714_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_714_inst
    process(iretire_state_reg_write_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_state_reg_write_710, R_one_1_713_wire_constant, tmp_var);
      EQ_u1_u1_714_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_723_inst flow-through 
    process(EQ_u1_u1_723_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_723_inst:flowthrough inputs: " & " iretire_state_reg_write_710 = "& Convert_SLV_To_Hex_String(iretire_state_reg_write_710) & " R_one_1_722_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_722_wire_constant) & " outputs:" & " EQ_u1_u1_723_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_723_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_723_inst
    process(iretire_state_reg_write_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_state_reg_write_710, R_one_1_722_wire_constant, tmp_var);
      EQ_u1_u1_723_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_732_inst flow-through 
    process(EQ_u1_u1_732_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_732_inst:flowthrough inputs: " & " iretire_state_reg_write_710 = "& Convert_SLV_To_Hex_String(iretire_state_reg_write_710) & " R_one_1_731_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_731_wire_constant) & " outputs:" & " EQ_u1_u1_732_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_732_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_732_inst
    process(iretire_state_reg_write_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_state_reg_write_710, R_one_1_731_wire_constant, tmp_var);
      EQ_u1_u1_732_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_741_inst flow-through 
    process(EQ_u1_u1_741_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_741_inst:flowthrough inputs: " & " iretire_state_reg_write_710 = "& Convert_SLV_To_Hex_String(iretire_state_reg_write_710) & " R_one_1_740_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_740_wire_constant) & " outputs:" & " EQ_u1_u1_741_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_741_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_741_inst
    process(iretire_state_reg_write_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_state_reg_write_710, R_one_1_740_wire_constant, tmp_var);
      EQ_u1_u1_741_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_762_inst flow-through 
    process(EQ_u1_u1_762_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_762_inst:flowthrough inputs: " & " iretire_state_reg_write_710 = "& Convert_SLV_To_Hex_String(iretire_state_reg_write_710) & " R_one_1_761_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_761_wire_constant) & " outputs:" & " EQ_u1_u1_762_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_762_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_762_inst
    process(iretire_state_reg_write_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_state_reg_write_710, R_one_1_761_wire_constant, tmp_var);
      EQ_u1_u1_762_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_771_inst flow-through 
    process(EQ_u1_u1_771_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_771_inst:flowthrough inputs: " & " iretire_state_reg_write_710 = "& Convert_SLV_To_Hex_String(iretire_state_reg_write_710) & " R_one_1_770_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_770_wire_constant) & " outputs:" & " EQ_u1_u1_771_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_771_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_771_inst
    process(iretire_state_reg_write_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_state_reg_write_710, R_one_1_770_wire_constant, tmp_var);
      EQ_u1_u1_771_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_803_inst flow-through 
    process(EQ_u1_u1_803_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_803_inst:flowthrough inputs: " & " is_Branch_538 = "& Convert_SLV_To_Hex_String(is_Branch_538) & " R_one_1_802_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_802_wire_constant) & " outputs:" & " EQ_u1_u1_803_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_803_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_803_inst
    process(is_Branch_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(is_Branch_538, R_one_1_802_wire_constant, tmp_var);
      EQ_u1_u1_803_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_806_inst flow-through 
    process(EQ_u1_u1_806_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_806_inst:flowthrough inputs: " & " ex_Unconditional_JUMP_buffer = "& Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_buffer) & " R_one_1_805_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_805_wire_constant) & " outputs:" & " EQ_u1_u1_806_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_806_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_806_inst
    process(ex_Unconditional_JUMP_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_Unconditional_JUMP_buffer, R_one_1_805_wire_constant, tmp_var);
      EQ_u1_u1_806_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_812_inst flow-through 
    process(EQ_u1_u1_812_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_812_inst:flowthrough inputs: " & " is_Branch_538 = "& Convert_SLV_To_Hex_String(is_Branch_538) & " R_one_1_811_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_811_wire_constant) & " outputs:" & " EQ_u1_u1_812_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_812_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_812_inst
    process(is_Branch_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(is_Branch_538, R_one_1_811_wire_constant, tmp_var);
      EQ_u1_u1_812_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_815_inst flow-through 
    process(EQ_u1_u1_815_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_815_inst:flowthrough inputs: " & " ex_Unconditional_JUMP_buffer = "& Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_buffer) & " R_one_1_814_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_814_wire_constant) & " outputs:" & " EQ_u1_u1_815_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_815_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_815_inst
    process(ex_Unconditional_JUMP_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_Unconditional_JUMP_buffer, R_one_1_814_wire_constant, tmp_var);
      EQ_u1_u1_815_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_821_inst flow-through 
    process(EQ_u1_u1_821_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_821_inst:flowthrough inputs: " & " is_Branch_538 = "& Convert_SLV_To_Hex_String(is_Branch_538) & " R_one_1_820_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_820_wire_constant) & " outputs:" & " EQ_u1_u1_821_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_821_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_821_inst
    process(is_Branch_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(is_Branch_538, R_one_1_820_wire_constant, tmp_var);
      EQ_u1_u1_821_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_824_inst flow-through 
    process(EQ_u1_u1_824_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_824_inst:flowthrough inputs: " & " ex_Unconditional_JUMP_buffer = "& Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_buffer) & " R_one_1_823_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_823_wire_constant) & " outputs:" & " EQ_u1_u1_824_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_824_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_824_inst
    process(ex_Unconditional_JUMP_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_Unconditional_JUMP_buffer, R_one_1_823_wire_constant, tmp_var);
      EQ_u1_u1_824_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_830_inst flow-through 
    process(EQ_u1_u1_830_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_830_inst:flowthrough inputs: " & " is_Branch_538 = "& Convert_SLV_To_Hex_String(is_Branch_538) & " R_one_1_829_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_829_wire_constant) & " outputs:" & " EQ_u1_u1_830_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_830_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_830_inst
    process(is_Branch_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(is_Branch_538, R_one_1_829_wire_constant, tmp_var);
      EQ_u1_u1_830_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_833_inst flow-through 
    process(EQ_u1_u1_833_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_833_inst:flowthrough inputs: " & " ex_Unconditional_JUMP_buffer = "& Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_buffer) & " R_one_1_832_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_832_wire_constant) & " outputs:" & " EQ_u1_u1_833_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_833_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_833_inst
    process(ex_Unconditional_JUMP_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_Unconditional_JUMP_buffer, R_one_1_832_wire_constant, tmp_var);
      EQ_u1_u1_833_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_839_inst flow-through 
    process(EQ_u1_u1_839_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_839_inst:flowthrough inputs: " & " is_Branch_538 = "& Convert_SLV_To_Hex_String(is_Branch_538) & " R_one_1_838_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_838_wire_constant) & " outputs:" & " EQ_u1_u1_839_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_839_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_839_inst
    process(is_Branch_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(is_Branch_538, R_one_1_838_wire_constant, tmp_var);
      EQ_u1_u1_839_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_842_inst flow-through 
    process(EQ_u1_u1_842_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_842_inst:flowthrough inputs: " & " ex_Unconditional_JUMP_buffer = "& Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_buffer) & " R_one_1_841_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_841_wire_constant) & " outputs:" & " EQ_u1_u1_842_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_842_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_842_inst
    process(ex_Unconditional_JUMP_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_Unconditional_JUMP_buffer, R_one_1_841_wire_constant, tmp_var);
      EQ_u1_u1_842_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_846_inst flow-through 
    process(EQ_u1_u1_846_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u1_u1_846_inst:flowthrough inputs: " & " stall_first_4_buffer = "& Convert_SLV_To_Hex_String(stall_first_4_buffer) & " R_one_1_845_wire_constant = "& Convert_SLV_To_Hex_String(R_one_1_845_wire_constant) & " outputs:" & " EQ_u1_u1_846_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_846_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_846_inst
    process(stall_first_4_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(stall_first_4_buffer, R_one_1_845_wire_constant, tmp_var);
      EQ_u1_u1_846_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_558_inst flow-through 
    process(EQ_u8_u1_558_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_558_inst:flowthrough inputs: " & " ex_opcode_542 = "& Convert_SLV_To_Hex_String(ex_opcode_542) & " R_CALL_557_wire_constant = "& Convert_SLV_To_Hex_String(R_CALL_557_wire_constant) & " outputs:" & " EQ_u8_u1_558_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_558_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_558_inst
    process(ex_opcode_542) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_opcode_542, R_CALL_557_wire_constant, tmp_var);
      EQ_u8_u1_558_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_561_inst flow-through 
    process(EQ_u8_u1_561_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_561_inst:flowthrough inputs: " & " ex_opcode_542 = "& Convert_SLV_To_Hex_String(ex_opcode_542) & " R_JMP_560_wire_constant = "& Convert_SLV_To_Hex_String(R_JMP_560_wire_constant) & " outputs:" & " EQ_u8_u1_561_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_561_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_561_inst
    process(ex_opcode_542) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_opcode_542, R_JMP_560_wire_constant, tmp_var);
      EQ_u8_u1_561_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_586_inst flow-through 
    process(EQ_u8_u1_586_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_586_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_SBIR_585_wire_constant = "& Convert_SLV_To_Hex_String(R_SBIR_585_wire_constant) & " outputs:" & " EQ_u8_u1_586_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_586_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_586_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_SBIR_585_wire_constant, tmp_var);
      EQ_u8_u1_586_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_589_inst flow-through 
    process(EQ_u8_u1_589_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_589_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_LOAD_588_wire_constant = "& Convert_SLV_To_Hex_String(R_LOAD_588_wire_constant) & " outputs:" & " EQ_u8_u1_589_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_589_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_589_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_LOAD_588_wire_constant, tmp_var);
      EQ_u8_u1_589_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_593_inst flow-through 
    process(EQ_u8_u1_593_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_593_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_L_AND_592_wire_constant = "& Convert_SLV_To_Hex_String(R_L_AND_592_wire_constant) & " outputs:" & " EQ_u8_u1_593_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_593_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_593_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_L_AND_592_wire_constant, tmp_var);
      EQ_u8_u1_593_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_597_inst flow-through 
    process(EQ_u8_u1_597_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_597_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_L_OR_596_wire_constant = "& Convert_SLV_To_Hex_String(R_L_OR_596_wire_constant) & " outputs:" & " EQ_u8_u1_597_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_597_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_597_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_L_OR_596_wire_constant, tmp_var);
      EQ_u8_u1_597_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_600_inst flow-through 
    process(EQ_u8_u1_600_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_600_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_L_XNOR_599_wire_constant = "& Convert_SLV_To_Hex_String(R_L_XNOR_599_wire_constant) & " outputs:" & " EQ_u8_u1_600_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_600_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_600_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_L_XNOR_599_wire_constant, tmp_var);
      EQ_u8_u1_600_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_604_inst flow-through 
    process(EQ_u8_u1_604_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_604_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_ADD_603_wire_constant = "& Convert_SLV_To_Hex_String(R_ADD_603_wire_constant) & " outputs:" & " EQ_u8_u1_604_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_604_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_604_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_ADD_603_wire_constant, tmp_var);
      EQ_u8_u1_604_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_609_inst flow-through 
    process(EQ_u8_u1_609_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_609_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_SUB_608_wire_constant = "& Convert_SLV_To_Hex_String(R_SUB_608_wire_constant) & " outputs:" & " EQ_u8_u1_609_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_609_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_609_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_SUB_608_wire_constant, tmp_var);
      EQ_u8_u1_609_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_612_inst flow-through 
    process(EQ_u8_u1_612_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_612_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_L_SLL_611_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SLL_611_wire_constant) & " outputs:" & " EQ_u8_u1_612_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_612_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_612_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_L_SLL_611_wire_constant, tmp_var);
      EQ_u8_u1_612_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_616_inst flow-through 
    process(EQ_u8_u1_616_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_616_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_L_SRL_615_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SRL_615_wire_constant) & " outputs:" & " EQ_u8_u1_616_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_616_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_616_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_L_SRL_615_wire_constant, tmp_var);
      EQ_u8_u1_616_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_620_inst flow-through 
    process(EQ_u8_u1_620_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_620_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_L_SRA_619_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SRA_619_wire_constant) & " outputs:" & " EQ_u8_u1_620_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_620_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_620_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_L_SRA_619_wire_constant, tmp_var);
      EQ_u8_u1_620_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_623_inst flow-through 
    process(EQ_u8_u1_623_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_623_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_CALL_622_wire_constant = "& Convert_SLV_To_Hex_String(R_CALL_622_wire_constant) & " outputs:" & " EQ_u8_u1_623_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_623_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_623_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_CALL_622_wire_constant, tmp_var);
      EQ_u8_u1_623_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_627_inst flow-through 
    process(EQ_u8_u1_627_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_627_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_CMP_626_wire_constant = "& Convert_SLV_To_Hex_String(R_CMP_626_wire_constant) & " outputs:" & " EQ_u8_u1_627_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_627_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_627_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_CMP_626_wire_constant, tmp_var);
      EQ_u8_u1_627_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_638_inst flow-through 
    process(EQ_u8_u1_638_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_638_inst:flowthrough inputs: " & " dcache_rd_582 = "& Convert_SLV_To_Hex_String(dcache_rd_582) & " ex_rs1_imm_546 = "& Convert_SLV_To_Hex_String(ex_rs1_imm_546) & " outputs:" & " EQ_u8_u1_638_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_638_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_638_inst
    process(dcache_rd_582, ex_rs1_imm_546) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_rd_582, ex_rs1_imm_546, tmp_var);
      EQ_u8_u1_638_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_647_inst flow-through 
    process(EQ_u8_u1_647_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_647_inst:flowthrough inputs: " & " dcache_rd_582 = "& Convert_SLV_To_Hex_String(dcache_rd_582) & " ex_rs2_550 = "& Convert_SLV_To_Hex_String(ex_rs2_550) & " outputs:" & " EQ_u8_u1_647_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_647_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_647_inst
    process(dcache_rd_582, ex_rs2_550) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_rd_582, ex_rs2_550, tmp_var);
      EQ_u8_u1_647_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_665_inst flow-through 
    process(EQ_u8_u1_665_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_665_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_SBIR_664_wire_constant = "& Convert_SLV_To_Hex_String(R_SBIR_664_wire_constant) & " outputs:" & " EQ_u8_u1_665_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_665_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_665_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_SBIR_664_wire_constant, tmp_var);
      EQ_u8_u1_665_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_668_inst flow-through 
    process(EQ_u8_u1_668_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_668_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_LOAD_667_wire_constant = "& Convert_SLV_To_Hex_String(R_LOAD_667_wire_constant) & " outputs:" & " EQ_u8_u1_668_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_668_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_668_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_LOAD_667_wire_constant, tmp_var);
      EQ_u8_u1_668_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_672_inst flow-through 
    process(EQ_u8_u1_672_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_672_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_L_AND_671_wire_constant = "& Convert_SLV_To_Hex_String(R_L_AND_671_wire_constant) & " outputs:" & " EQ_u8_u1_672_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_672_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_672_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_L_AND_671_wire_constant, tmp_var);
      EQ_u8_u1_672_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_676_inst flow-through 
    process(EQ_u8_u1_676_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_676_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_L_OR_675_wire_constant = "& Convert_SLV_To_Hex_String(R_L_OR_675_wire_constant) & " outputs:" & " EQ_u8_u1_676_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_676_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_676_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_L_OR_675_wire_constant, tmp_var);
      EQ_u8_u1_676_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_679_inst flow-through 
    process(EQ_u8_u1_679_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_679_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_L_XNOR_678_wire_constant = "& Convert_SLV_To_Hex_String(R_L_XNOR_678_wire_constant) & " outputs:" & " EQ_u8_u1_679_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_679_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_679_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_L_XNOR_678_wire_constant, tmp_var);
      EQ_u8_u1_679_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_683_inst flow-through 
    process(EQ_u8_u1_683_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_683_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_ADD_682_wire_constant = "& Convert_SLV_To_Hex_String(R_ADD_682_wire_constant) & " outputs:" & " EQ_u8_u1_683_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_683_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_683_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_ADD_682_wire_constant, tmp_var);
      EQ_u8_u1_683_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_688_inst flow-through 
    process(EQ_u8_u1_688_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_688_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_SUB_687_wire_constant = "& Convert_SLV_To_Hex_String(R_SUB_687_wire_constant) & " outputs:" & " EQ_u8_u1_688_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_688_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_688_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_SUB_687_wire_constant, tmp_var);
      EQ_u8_u1_688_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_691_inst flow-through 
    process(EQ_u8_u1_691_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_691_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_L_SLL_690_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SLL_690_wire_constant) & " outputs:" & " EQ_u8_u1_691_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_691_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_691_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_L_SLL_690_wire_constant, tmp_var);
      EQ_u8_u1_691_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_695_inst flow-through 
    process(EQ_u8_u1_695_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_695_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_L_SRL_694_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SRL_694_wire_constant) & " outputs:" & " EQ_u8_u1_695_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_695_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_695_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_L_SRL_694_wire_constant, tmp_var);
      EQ_u8_u1_695_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_699_inst flow-through 
    process(EQ_u8_u1_699_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_699_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_L_SRA_698_wire_constant = "& Convert_SLV_To_Hex_String(R_L_SRA_698_wire_constant) & " outputs:" & " EQ_u8_u1_699_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_699_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_699_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_L_SRA_698_wire_constant, tmp_var);
      EQ_u8_u1_699_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_702_inst flow-through 
    process(EQ_u8_u1_702_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_702_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_CALL_701_wire_constant = "& Convert_SLV_To_Hex_String(R_CALL_701_wire_constant) & " outputs:" & " EQ_u8_u1_702_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_702_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_702_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_CALL_701_wire_constant, tmp_var);
      EQ_u8_u1_702_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_706_inst flow-through 
    process(EQ_u8_u1_706_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_706_inst:flowthrough inputs: " & " iretire_opcode_653 = "& Convert_SLV_To_Hex_String(iretire_opcode_653) & " R_CMP_705_wire_constant = "& Convert_SLV_To_Hex_String(R_CMP_705_wire_constant) & " outputs:" & " EQ_u8_u1_706_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_706_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_706_inst
    process(iretire_opcode_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_opcode_653, R_CMP_705_wire_constant, tmp_var);
      EQ_u8_u1_706_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_717_inst flow-through 
    process(EQ_u8_u1_717_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_717_inst:flowthrough inputs: " & " iretire_rd_661 = "& Convert_SLV_To_Hex_String(iretire_rd_661) & " ex_rs1_imm_546 = "& Convert_SLV_To_Hex_String(ex_rs1_imm_546) & " outputs:" & " EQ_u8_u1_717_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_717_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_717_inst
    process(iretire_rd_661, ex_rs1_imm_546) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_rd_661, ex_rs1_imm_546, tmp_var);
      EQ_u8_u1_717_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_726_inst flow-through 
    process(EQ_u8_u1_726_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_726_inst:flowthrough inputs: " & " iretire_rd_661 = "& Convert_SLV_To_Hex_String(iretire_rd_661) & " ex_rs2_550 = "& Convert_SLV_To_Hex_String(ex_rs2_550) & " outputs:" & " EQ_u8_u1_726_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_726_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_726_inst
    process(iretire_rd_661, ex_rs2_550) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_rd_661, ex_rs2_550, tmp_var);
      EQ_u8_u1_726_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_735_inst flow-through 
    process(EQ_u8_u1_735_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_735_inst:flowthrough inputs: " & " dcache_rs1_imm_574 = "& Convert_SLV_To_Hex_String(dcache_rs1_imm_574) & " iretire_rd_661 = "& Convert_SLV_To_Hex_String(iretire_rd_661) & " outputs:" & " EQ_u8_u1_735_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_735_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_735_inst
    process(dcache_rs1_imm_574, iretire_rd_661) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_rs1_imm_574, iretire_rd_661, tmp_var);
      EQ_u8_u1_735_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_744_inst flow-through 
    process(EQ_u8_u1_744_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_744_inst:flowthrough inputs: " & " dcache_rs2_578 = "& Convert_SLV_To_Hex_String(dcache_rs2_578) & " iretire_rd_661 = "& Convert_SLV_To_Hex_String(iretire_rd_661) & " outputs:" & " EQ_u8_u1_744_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_744_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_744_inst
    process(dcache_rs2_578, iretire_rd_661) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_rs2_578, iretire_rd_661, tmp_var);
      EQ_u8_u1_744_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_765_inst flow-through 
    process(EQ_u8_u1_765_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_765_inst:flowthrough inputs: " & " iretire_rd_661 = "& Convert_SLV_To_Hex_String(iretire_rd_661) & " iregfile_rs1_imm_754 = "& Convert_SLV_To_Hex_String(iregfile_rs1_imm_754) & " outputs:" & " EQ_u8_u1_765_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_765_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_765_inst
    process(iretire_rd_661, iregfile_rs1_imm_754) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_rd_661, iregfile_rs1_imm_754, tmp_var);
      EQ_u8_u1_765_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_774_inst flow-through 
    process(EQ_u8_u1_774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_774_inst:flowthrough inputs: " & " iretire_rd_661 = "& Convert_SLV_To_Hex_String(iretire_rd_661) & " iregfile_rs2_758 = "& Convert_SLV_To_Hex_String(iregfile_rs2_758) & " outputs:" & " EQ_u8_u1_774_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_774_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_774_inst
    process(iretire_rd_661, iregfile_rs2_758) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_rd_661, iregfile_rs2_758, tmp_var);
      EQ_u8_u1_774_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_780_inst flow-through 
    process(EQ_u8_u1_780_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_780_inst:flowthrough inputs: " & " ex_opcode_542 = "& Convert_SLV_To_Hex_String(ex_opcode_542) & " R_LOAD_779_wire_constant = "& Convert_SLV_To_Hex_String(R_LOAD_779_wire_constant) & " outputs:" & " EQ_u8_u1_780_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_780_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_780_inst
    process(ex_opcode_542) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ex_opcode_542, R_LOAD_779_wire_constant, tmp_var);
      EQ_u8_u1_780_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_783_inst flow-through 
    process(EQ_u8_u1_783_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_783_inst:flowthrough inputs: " & " iregfile_opcode_750 = "& Convert_SLV_To_Hex_String(iregfile_opcode_750) & " R_zero_8_782_wire_constant = "& Convert_SLV_To_Hex_String(R_zero_8_782_wire_constant) & " outputs:" & " EQ_u8_u1_783_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_783_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_783_inst
    process(iregfile_opcode_750) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iregfile_opcode_750, R_zero_8_782_wire_constant, tmp_var);
      EQ_u8_u1_783_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_788_inst flow-through 
    process(EQ_u8_u1_788_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_788_inst:flowthrough inputs: " & " iregfile_opcode_750 = "& Convert_SLV_To_Hex_String(iregfile_opcode_750) & " R_STORE_787_wire_constant = "& Convert_SLV_To_Hex_String(R_STORE_787_wire_constant) & " outputs:" & " EQ_u8_u1_788_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_788_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_788_inst
    process(iregfile_opcode_750) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iregfile_opcode_750, R_STORE_787_wire_constant, tmp_var);
      EQ_u8_u1_788_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_792_inst flow-through 
    process(EQ_u8_u1_792_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_792_inst:flowthrough inputs: " & " iretire_rs1_imm_657 = "& Convert_SLV_To_Hex_String(iretire_rs1_imm_657) & " ex_rd_554 = "& Convert_SLV_To_Hex_String(ex_rd_554) & " outputs:" & " EQ_u8_u1_792_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_792_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_792_inst
    process(iretire_rs1_imm_657, ex_rd_554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iretire_rs1_imm_657, ex_rd_554, tmp_var);
      EQ_u8_u1_792_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_795_inst flow-through 
    process(EQ_u8_u1_795_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_795_inst:flowthrough inputs: " & " iregfile_rs2_758 = "& Convert_SLV_To_Hex_String(iregfile_rs2_758) & " ex_rd_554 = "& Convert_SLV_To_Hex_String(ex_rd_554) & " outputs:" & " EQ_u8_u1_795_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_795_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_795_inst
    process(iregfile_rs2_758, ex_rd_554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iregfile_rs2_758, ex_rd_554, tmp_var);
      EQ_u8_u1_795_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_868_inst flow-through 
    process(EQ_u8_u1_868_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_868_inst:flowthrough inputs: " & " iregfile_state_opcode_864 = "& Convert_SLV_To_Hex_String(iregfile_state_opcode_864) & " konst_867_wire_constant = "& Convert_SLV_To_Hex_String(konst_867_wire_constant) & " outputs:" & " EQ_u8_u1_868_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_868_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_868_inst
    process(iregfile_state_opcode_864) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iregfile_state_opcode_864, konst_867_wire_constant, tmp_var);
      EQ_u8_u1_868_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_876_inst flow-through 
    process(EQ_u8_u1_876_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_876_inst:flowthrough inputs: " & " iregfile_state_opcode_864 = "& Convert_SLV_To_Hex_String(iregfile_state_opcode_864) & " konst_875_wire_constant = "& Convert_SLV_To_Hex_String(konst_875_wire_constant) & " outputs:" & " EQ_u8_u1_876_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_876_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_876_inst
    process(iregfile_state_opcode_864) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iregfile_state_opcode_864, konst_875_wire_constant, tmp_var);
      EQ_u8_u1_876_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_907_inst flow-through 
    process(EQ_u8_u1_907_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:EQ_u8_u1_907_inst:flowthrough inputs: " & " dcache_opcode_570 = "& Convert_SLV_To_Hex_String(dcache_opcode_570) & " R_STORE_906_wire_constant = "& Convert_SLV_To_Hex_String(R_STORE_906_wire_constant) & " outputs:" & " EQ_u8_u1_907_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_907_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_907_inst
    process(dcache_opcode_570) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dcache_opcode_570, R_STORE_906_wire_constant, tmp_var);
      EQ_u8_u1_907_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_784_inst flow-through 
    process(NOT_u1_u1_784_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:NOT_u1_u1_784_inst:flowthrough inputs: " & " EQ_u8_u1_783_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_783_wire) & " outputs:" & " NOT_u1_u1_784_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_784_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_784_inst
    process(EQ_u8_u1_783_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", EQ_u8_u1_783_wire, tmp_var);
      NOT_u1_u1_784_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator NOT_u1_u1_789_inst flow-through 
    process(NOT_u1_u1_789_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:NOT_u1_u1_789_inst:flowthrough inputs: " & " EQ_u8_u1_788_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_788_wire) & " outputs:" & " NOT_u1_u1_789_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_789_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_789_inst
    process(EQ_u8_u1_788_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", EQ_u8_u1_788_wire, tmp_var);
      NOT_u1_u1_789_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator OR_u1_u1_562_inst flow-through 
    process(ex_Unconditional_JUMP_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_562_inst:flowthrough inputs: " & " EQ_u8_u1_558_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_558_wire) & " EQ_u8_u1_561_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_561_wire) & " outputs:" & " ex_Unconditional_JUMP_buffer= "  & Convert_SLV_To_Hex_String(ex_Unconditional_JUMP_buffer));
      --
    end process; 
    -- binary operator OR_u1_u1_562_inst
    process(EQ_u8_u1_558_wire, EQ_u8_u1_561_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_558_wire, EQ_u8_u1_561_wire, tmp_var);
      ex_Unconditional_JUMP_buffer <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_590_inst flow-through 
    process(OR_u1_u1_590_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_590_inst:flowthrough inputs: " & " EQ_u8_u1_586_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_586_wire) & " EQ_u8_u1_589_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_589_wire) & " outputs:" & " OR_u1_u1_590_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_590_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_590_inst
    process(EQ_u8_u1_586_wire, EQ_u8_u1_589_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_586_wire, EQ_u8_u1_589_wire, tmp_var);
      OR_u1_u1_590_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_594_inst flow-through 
    process(OR_u1_u1_594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_594_inst:flowthrough inputs: " & " OR_u1_u1_590_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_590_wire) & " EQ_u8_u1_593_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_593_wire) & " outputs:" & " OR_u1_u1_594_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_594_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_594_inst
    process(OR_u1_u1_590_wire, EQ_u8_u1_593_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_590_wire, EQ_u8_u1_593_wire, tmp_var);
      OR_u1_u1_594_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_601_inst flow-through 
    process(OR_u1_u1_601_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_601_inst:flowthrough inputs: " & " EQ_u8_u1_597_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_597_wire) & " EQ_u8_u1_600_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_600_wire) & " outputs:" & " OR_u1_u1_601_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_601_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_601_inst
    process(EQ_u8_u1_597_wire, EQ_u8_u1_600_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_597_wire, EQ_u8_u1_600_wire, tmp_var);
      OR_u1_u1_601_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_605_inst flow-through 
    process(OR_u1_u1_605_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_605_inst:flowthrough inputs: " & " OR_u1_u1_601_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_601_wire) & " EQ_u8_u1_604_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_604_wire) & " outputs:" & " OR_u1_u1_605_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_605_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_605_inst
    process(OR_u1_u1_601_wire, EQ_u8_u1_604_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_601_wire, EQ_u8_u1_604_wire, tmp_var);
      OR_u1_u1_605_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_606_inst flow-through 
    process(OR_u1_u1_606_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_606_inst:flowthrough inputs: " & " OR_u1_u1_594_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_594_wire) & " OR_u1_u1_605_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_605_wire) & " outputs:" & " OR_u1_u1_606_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_606_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_606_inst
    process(OR_u1_u1_594_wire, OR_u1_u1_605_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_594_wire, OR_u1_u1_605_wire, tmp_var);
      OR_u1_u1_606_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_613_inst flow-through 
    process(OR_u1_u1_613_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_613_inst:flowthrough inputs: " & " EQ_u8_u1_609_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_609_wire) & " EQ_u8_u1_612_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_612_wire) & " outputs:" & " OR_u1_u1_613_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_613_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_613_inst
    process(EQ_u8_u1_609_wire, EQ_u8_u1_612_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_609_wire, EQ_u8_u1_612_wire, tmp_var);
      OR_u1_u1_613_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_617_inst flow-through 
    process(OR_u1_u1_617_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_617_inst:flowthrough inputs: " & " OR_u1_u1_613_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_613_wire) & " EQ_u8_u1_616_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_616_wire) & " outputs:" & " OR_u1_u1_617_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_617_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_617_inst
    process(OR_u1_u1_613_wire, EQ_u8_u1_616_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_613_wire, EQ_u8_u1_616_wire, tmp_var);
      OR_u1_u1_617_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_624_inst flow-through 
    process(OR_u1_u1_624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_624_inst:flowthrough inputs: " & " EQ_u8_u1_620_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_620_wire) & " EQ_u8_u1_623_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_623_wire) & " outputs:" & " OR_u1_u1_624_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_624_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_624_inst
    process(EQ_u8_u1_620_wire, EQ_u8_u1_623_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_620_wire, EQ_u8_u1_623_wire, tmp_var);
      OR_u1_u1_624_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_628_inst flow-through 
    process(OR_u1_u1_628_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_628_inst:flowthrough inputs: " & " OR_u1_u1_624_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_624_wire) & " EQ_u8_u1_627_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_627_wire) & " outputs:" & " OR_u1_u1_628_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_628_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_628_inst
    process(OR_u1_u1_624_wire, EQ_u8_u1_627_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_624_wire, EQ_u8_u1_627_wire, tmp_var);
      OR_u1_u1_628_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_629_inst flow-through 
    process(OR_u1_u1_629_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_629_inst:flowthrough inputs: " & " OR_u1_u1_617_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_617_wire) & " OR_u1_u1_628_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_628_wire) & " outputs:" & " OR_u1_u1_629_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_629_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_629_inst
    process(OR_u1_u1_617_wire, OR_u1_u1_628_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_617_wire, OR_u1_u1_628_wire, tmp_var);
      OR_u1_u1_629_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_630_inst flow-through 
    process(dcache_state_reg_write_631) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_630_inst:flowthrough inputs: " & " OR_u1_u1_606_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_606_wire) & " OR_u1_u1_629_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_629_wire) & " outputs:" & " dcache_state_reg_write_631= "  & Convert_SLV_To_Hex_String(dcache_state_reg_write_631));
      --
    end process; 
    -- binary operator OR_u1_u1_630_inst
    process(OR_u1_u1_606_wire, OR_u1_u1_629_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_606_wire, OR_u1_u1_629_wire, tmp_var);
      dcache_state_reg_write_631 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_669_inst flow-through 
    process(OR_u1_u1_669_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_669_inst:flowthrough inputs: " & " EQ_u8_u1_665_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_665_wire) & " EQ_u8_u1_668_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_668_wire) & " outputs:" & " OR_u1_u1_669_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_669_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_669_inst
    process(EQ_u8_u1_665_wire, EQ_u8_u1_668_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_665_wire, EQ_u8_u1_668_wire, tmp_var);
      OR_u1_u1_669_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_673_inst flow-through 
    process(OR_u1_u1_673_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_673_inst:flowthrough inputs: " & " OR_u1_u1_669_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_669_wire) & " EQ_u8_u1_672_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_672_wire) & " outputs:" & " OR_u1_u1_673_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_673_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_673_inst
    process(OR_u1_u1_669_wire, EQ_u8_u1_672_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_669_wire, EQ_u8_u1_672_wire, tmp_var);
      OR_u1_u1_673_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_680_inst flow-through 
    process(OR_u1_u1_680_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_680_inst:flowthrough inputs: " & " EQ_u8_u1_676_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_676_wire) & " EQ_u8_u1_679_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_679_wire) & " outputs:" & " OR_u1_u1_680_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_680_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_680_inst
    process(EQ_u8_u1_676_wire, EQ_u8_u1_679_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_676_wire, EQ_u8_u1_679_wire, tmp_var);
      OR_u1_u1_680_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_684_inst flow-through 
    process(OR_u1_u1_684_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_684_inst:flowthrough inputs: " & " OR_u1_u1_680_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_680_wire) & " EQ_u8_u1_683_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_683_wire) & " outputs:" & " OR_u1_u1_684_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_684_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_684_inst
    process(OR_u1_u1_680_wire, EQ_u8_u1_683_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_680_wire, EQ_u8_u1_683_wire, tmp_var);
      OR_u1_u1_684_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_685_inst flow-through 
    process(OR_u1_u1_685_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_685_inst:flowthrough inputs: " & " OR_u1_u1_673_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_673_wire) & " OR_u1_u1_684_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_684_wire) & " outputs:" & " OR_u1_u1_685_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_685_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_685_inst
    process(OR_u1_u1_673_wire, OR_u1_u1_684_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_673_wire, OR_u1_u1_684_wire, tmp_var);
      OR_u1_u1_685_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_692_inst flow-through 
    process(OR_u1_u1_692_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_692_inst:flowthrough inputs: " & " EQ_u8_u1_688_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_688_wire) & " EQ_u8_u1_691_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_691_wire) & " outputs:" & " OR_u1_u1_692_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_692_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_692_inst
    process(EQ_u8_u1_688_wire, EQ_u8_u1_691_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_688_wire, EQ_u8_u1_691_wire, tmp_var);
      OR_u1_u1_692_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_696_inst flow-through 
    process(OR_u1_u1_696_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_696_inst:flowthrough inputs: " & " OR_u1_u1_692_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_692_wire) & " EQ_u8_u1_695_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_695_wire) & " outputs:" & " OR_u1_u1_696_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_696_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_696_inst
    process(OR_u1_u1_692_wire, EQ_u8_u1_695_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_692_wire, EQ_u8_u1_695_wire, tmp_var);
      OR_u1_u1_696_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_703_inst flow-through 
    process(OR_u1_u1_703_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_703_inst:flowthrough inputs: " & " EQ_u8_u1_699_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_699_wire) & " EQ_u8_u1_702_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_702_wire) & " outputs:" & " OR_u1_u1_703_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_703_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_703_inst
    process(EQ_u8_u1_699_wire, EQ_u8_u1_702_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_699_wire, EQ_u8_u1_702_wire, tmp_var);
      OR_u1_u1_703_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_707_inst flow-through 
    process(OR_u1_u1_707_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_707_inst:flowthrough inputs: " & " OR_u1_u1_703_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_703_wire) & " EQ_u8_u1_706_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_706_wire) & " outputs:" & " OR_u1_u1_707_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_707_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_707_inst
    process(OR_u1_u1_703_wire, EQ_u8_u1_706_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_703_wire, EQ_u8_u1_706_wire, tmp_var);
      OR_u1_u1_707_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_708_inst flow-through 
    process(OR_u1_u1_708_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_708_inst:flowthrough inputs: " & " OR_u1_u1_696_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_696_wire) & " OR_u1_u1_707_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_707_wire) & " outputs:" & " OR_u1_u1_708_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_708_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_708_inst
    process(OR_u1_u1_696_wire, OR_u1_u1_707_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_696_wire, OR_u1_u1_707_wire, tmp_var);
      OR_u1_u1_708_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_709_inst flow-through 
    process(iretire_state_reg_write_710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_709_inst:flowthrough inputs: " & " OR_u1_u1_685_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_685_wire) & " OR_u1_u1_708_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_708_wire) & " outputs:" & " iretire_state_reg_write_710= "  & Convert_SLV_To_Hex_String(iretire_state_reg_write_710));
      --
    end process; 
    -- binary operator OR_u1_u1_709_inst
    process(OR_u1_u1_685_wire, OR_u1_u1_708_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_685_wire, OR_u1_u1_708_wire, tmp_var);
      iretire_state_reg_write_710 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_796_inst flow-through 
    process(OR_u1_u1_796_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_796_inst:flowthrough inputs: " & " EQ_u8_u1_792_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_792_wire) & " EQ_u8_u1_795_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_795_wire) & " outputs:" & " OR_u1_u1_796_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_796_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_796_inst
    process(EQ_u8_u1_792_wire, EQ_u8_u1_795_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_792_wire, EQ_u8_u1_795_wire, tmp_var);
      OR_u1_u1_796_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_807_inst flow-through 
    process(flush_ifetch_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_807_inst:flowthrough inputs: " & " EQ_u1_u1_803_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_803_wire) & " EQ_u1_u1_806_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_806_wire) & " outputs:" & " flush_ifetch_buffer= "  & Convert_SLV_To_Hex_String(flush_ifetch_buffer));
      --
    end process; 
    -- binary operator OR_u1_u1_807_inst
    process(EQ_u1_u1_803_wire, EQ_u1_u1_806_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u1_u1_803_wire, EQ_u1_u1_806_wire, tmp_var);
      flush_ifetch_buffer <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_816_inst flow-through 
    process(flush_icache_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_816_inst:flowthrough inputs: " & " EQ_u1_u1_812_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_812_wire) & " EQ_u1_u1_815_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_815_wire) & " outputs:" & " flush_icache_buffer= "  & Convert_SLV_To_Hex_String(flush_icache_buffer));
      --
    end process; 
    -- binary operator OR_u1_u1_816_inst
    process(EQ_u1_u1_812_wire, EQ_u1_u1_815_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u1_u1_812_wire, EQ_u1_u1_815_wire, tmp_var);
      flush_icache_buffer <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_825_inst flow-through 
    process(flush_idecode_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_825_inst:flowthrough inputs: " & " EQ_u1_u1_821_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_821_wire) & " EQ_u1_u1_824_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_824_wire) & " outputs:" & " flush_idecode_buffer= "  & Convert_SLV_To_Hex_String(flush_idecode_buffer));
      --
    end process; 
    -- binary operator OR_u1_u1_825_inst
    process(EQ_u1_u1_821_wire, EQ_u1_u1_824_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u1_u1_821_wire, EQ_u1_u1_824_wire, tmp_var);
      flush_idecode_buffer <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_834_inst flow-through 
    process(flush_reg_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_834_inst:flowthrough inputs: " & " EQ_u1_u1_830_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_830_wire) & " EQ_u1_u1_833_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_833_wire) & " outputs:" & " flush_reg_buffer= "  & Convert_SLV_To_Hex_String(flush_reg_buffer));
      --
    end process; 
    -- binary operator OR_u1_u1_834_inst
    process(EQ_u1_u1_830_wire, EQ_u1_u1_833_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u1_u1_830_wire, EQ_u1_u1_833_wire, tmp_var);
      flush_reg_buffer <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_843_inst flow-through 
    process(OR_u1_u1_843_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_843_inst:flowthrough inputs: " & " EQ_u1_u1_839_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_839_wire) & " EQ_u1_u1_842_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_842_wire) & " outputs:" & " OR_u1_u1_843_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_843_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_843_inst
    process(EQ_u1_u1_839_wire, EQ_u1_u1_842_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u1_u1_839_wire, EQ_u1_u1_842_wire, tmp_var);
      OR_u1_u1_843_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_847_inst flow-through 
    process(flush_iexec_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:scoreBoard:DP:OR_u1_u1_847_inst:flowthrough inputs: " & " OR_u1_u1_843_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_843_wire) & " EQ_u1_u1_846_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_846_wire) & " outputs:" & " flush_iexec_buffer= "  & Convert_SLV_To_Hex_String(flush_iexec_buffer));
      --
    end process; 
    -- binary operator OR_u1_u1_847_inst
    process(OR_u1_u1_843_wire, EQ_u1_u1_846_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_843_wire, EQ_u1_u1_846_wire, tmp_var);
      flush_iexec_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end scoreBoard_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    accessMem_request_pipe_write_data: in std_logic_vector(63 downto 0);
    accessMem_request_pipe_write_req : in std_logic_vector(0 downto 0);
    accessMem_request_pipe_write_ack : out std_logic_vector(0 downto 0);
    accessMem_response_pipe_read_data: out std_logic_vector(31 downto 0);
    accessMem_response_pipe_read_req : in std_logic_vector(0 downto 0);
    accessMem_response_pipe_read_ack : out std_logic_vector(0 downto 0);
    accessReg_request_pipe_write_data: in std_logic_vector(63 downto 0);
    accessReg_request_pipe_write_req : in std_logic_vector(0 downto 0);
    accessReg_request_pipe_write_ack : out std_logic_vector(0 downto 0);
    accessReg_response1_pipe_read_data: out std_logic_vector(31 downto 0);
    accessReg_response1_pipe_read_req : in std_logic_vector(0 downto 0);
    accessReg_response1_pipe_read_ack : out std_logic_vector(0 downto 0);
    accessReg_response2_pipe_read_data: out std_logic_vector(31 downto 0);
    accessReg_response2_pipe_read_req : in std_logic_vector(0 downto 0);
    accessReg_response2_pipe_read_ack : out std_logic_vector(0 downto 0);
    processor_result_pipe_read_data: out std_logic_vector(31 downto 0);
    processor_result_pipe_read_req : in std_logic_vector(0 downto 0);
    processor_result_pipe_read_ack : out std_logic_vector(0 downto 0);
    start_processor_pipe_write_data: in std_logic_vector(7 downto 0);
    start_processor_pipe_write_req : in std_logic_vector(0 downto 0);
    start_processor_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(5 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(5 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module accessMem
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(9 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMem
  signal accessMem_read_write_bar :  std_logic_vector(0 downto 0);
  signal accessMem_addr :  std_logic_vector(9 downto 0);
  signal accessMem_write_data :  std_logic_vector(31 downto 0);
  signal accessMem_read_data :  std_logic_vector(31 downto 0);
  signal accessMem_in_args    : std_logic_vector(42 downto 0);
  signal accessMem_out_args   : std_logic_vector(31 downto 0);
  signal accessMem_tag_in    : std_logic_vector(3 downto 0) := (others => '0');
  signal accessMem_tag_out   : std_logic_vector(3 downto 0);
  signal accessMem_start_req : std_logic;
  signal accessMem_start_ack : std_logic;
  signal accessMem_fin_req   : std_logic;
  signal accessMem_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMem
  signal accessMem_call_reqs: std_logic_vector(1 downto 0);
  signal accessMem_call_acks: std_logic_vector(1 downto 0);
  signal accessMem_return_reqs: std_logic_vector(1 downto 0);
  signal accessMem_return_acks: std_logic_vector(1 downto 0);
  signal accessMem_call_data: std_logic_vector(85 downto 0);
  signal accessMem_call_tag: std_logic_vector(3 downto 0);
  signal accessMem_return_data: std_logic_vector(63 downto 0);
  signal accessMem_return_tag: std_logic_vector(3 downto 0);
  -- declarations related to module accessReg
  component accessReg is -- 
    generic (tag_length : integer); 
    port ( -- 
      valid_1 : in  std_logic_vector(0 downto 0);
      addr_1 : in  std_logic_vector(7 downto 0);
      valid_2 : in  std_logic_vector(0 downto 0);
      addr_2 : in  std_logic_vector(7 downto 0);
      valid_w : in  std_logic_vector(0 downto 0);
      addr_w : in  std_logic_vector(7 downto 0);
      data_to_be_written : in  std_logic_vector(31 downto 0);
      read_data_1 : out  std_logic_vector(31 downto 0);
      read_data_2 : out  std_logic_vector(31 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessReg
  signal accessReg_valid_1 :  std_logic_vector(0 downto 0);
  signal accessReg_addr_1 :  std_logic_vector(7 downto 0);
  signal accessReg_valid_2 :  std_logic_vector(0 downto 0);
  signal accessReg_addr_2 :  std_logic_vector(7 downto 0);
  signal accessReg_valid_w :  std_logic_vector(0 downto 0);
  signal accessReg_addr_w :  std_logic_vector(7 downto 0);
  signal accessReg_data_to_be_written :  std_logic_vector(31 downto 0);
  signal accessReg_read_data_1 :  std_logic_vector(31 downto 0);
  signal accessReg_read_data_2 :  std_logic_vector(31 downto 0);
  signal accessReg_in_args    : std_logic_vector(58 downto 0);
  signal accessReg_out_args   : std_logic_vector(63 downto 0);
  signal accessReg_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessReg_tag_out   : std_logic_vector(2 downto 0);
  signal accessReg_start_req : std_logic;
  signal accessReg_start_ack : std_logic;
  signal accessReg_fin_req   : std_logic;
  signal accessReg_fin_ack : std_logic;
  -- caller side aggregated signals for module accessReg
  signal accessReg_call_reqs: std_logic_vector(1 downto 0);
  signal accessReg_call_acks: std_logic_vector(1 downto 0);
  signal accessReg_return_reqs: std_logic_vector(1 downto 0);
  signal accessReg_return_acks: std_logic_vector(1 downto 0);
  signal accessReg_call_data: std_logic_vector(117 downto 0);
  signal accessReg_call_tag: std_logic_vector(1 downto 0);
  signal accessReg_return_data: std_logic_vector(127 downto 0);
  signal accessReg_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module iExecStage
  component iExecStage is -- 
    generic (tag_length : integer); 
    port ( -- 
      iexec_state : in  std_logic_vector(105 downto 0);
      iexec_rd1_final : in  std_logic_vector(31 downto 0);
      iexec_rd2_final : in  std_logic_vector(31 downto 0);
      next_dcache_state : out  std_logic_vector(138 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module iExecStage
  signal iExecStage_iexec_state :  std_logic_vector(105 downto 0);
  signal iExecStage_iexec_rd1_final :  std_logic_vector(31 downto 0);
  signal iExecStage_iexec_rd2_final :  std_logic_vector(31 downto 0);
  signal iExecStage_next_dcache_state :  std_logic_vector(138 downto 0);
  signal iExecStage_in_args    : std_logic_vector(169 downto 0);
  signal iExecStage_out_args   : std_logic_vector(138 downto 0);
  signal iExecStage_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal iExecStage_tag_out   : std_logic_vector(1 downto 0);
  signal iExecStage_start_req : std_logic;
  signal iExecStage_start_ack : std_logic;
  signal iExecStage_fin_req   : std_logic;
  signal iExecStage_fin_ack : std_logic;
  -- caller side aggregated signals for module iExecStage
  signal iExecStage_call_reqs: std_logic_vector(0 downto 0);
  signal iExecStage_call_acks: std_logic_vector(0 downto 0);
  signal iExecStage_return_reqs: std_logic_vector(0 downto 0);
  signal iExecStage_return_acks: std_logic_vector(0 downto 0);
  signal iExecStage_call_data: std_logic_vector(169 downto 0);
  signal iExecStage_call_tag: std_logic_vector(0 downto 0);
  signal iExecStage_return_data: std_logic_vector(138 downto 0);
  signal iExecStage_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module memAccessDaemon
  component memAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      accessMem_request_pipe_read_req : out  std_logic_vector(0 downto 0);
      accessMem_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
      accessMem_request_pipe_read_data : in   std_logic_vector(63 downto 0);
      accessMem_response_pipe_write_req : out  std_logic_vector(0 downto 0);
      accessMem_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
      accessMem_response_pipe_write_data : out  std_logic_vector(31 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(42 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(31 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module memAccessDaemon
  signal memAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal memAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal memAccessDaemon_start_req : std_logic;
  signal memAccessDaemon_start_ack : std_logic;
  signal memAccessDaemon_fin_req   : std_logic;
  signal memAccessDaemon_fin_ack : std_logic;
  -- declarations related to module processor_daemon
  component processor_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_processor_pipe_read_req : out  std_logic_vector(0 downto 0);
      start_processor_pipe_read_ack : in   std_logic_vector(0 downto 0);
      start_processor_pipe_read_data : in   std_logic_vector(7 downto 0);
      processor_result_pipe_write_req : out  std_logic_vector(0 downto 0);
      processor_result_pipe_write_ack : in   std_logic_vector(0 downto 0);
      processor_result_pipe_write_data : out  std_logic_vector(31 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(42 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(31 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      iExecStage_call_reqs : out  std_logic_vector(0 downto 0);
      iExecStage_call_acks : in   std_logic_vector(0 downto 0);
      iExecStage_call_data : out  std_logic_vector(169 downto 0);
      iExecStage_call_tag  :  out  std_logic_vector(0 downto 0);
      iExecStage_return_reqs : out  std_logic_vector(0 downto 0);
      iExecStage_return_acks : in   std_logic_vector(0 downto 0);
      iExecStage_return_data : in   std_logic_vector(138 downto 0);
      iExecStage_return_tag :  in   std_logic_vector(0 downto 0);
      accessReg_call_reqs : out  std_logic_vector(0 downto 0);
      accessReg_call_acks : in   std_logic_vector(0 downto 0);
      accessReg_call_data : out  std_logic_vector(58 downto 0);
      accessReg_call_tag  :  out  std_logic_vector(0 downto 0);
      accessReg_return_reqs : out  std_logic_vector(0 downto 0);
      accessReg_return_acks : in   std_logic_vector(0 downto 0);
      accessReg_return_data : in   std_logic_vector(63 downto 0);
      accessReg_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module processor_daemon
  signal processor_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal processor_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal processor_daemon_start_req : std_logic;
  signal processor_daemon_start_ack : std_logic;
  signal processor_daemon_fin_req   : std_logic;
  signal processor_daemon_fin_ack : std_logic;
  -- declarations related to module regAccessDaemon
  component regAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      accessReg_request_pipe_read_req : out  std_logic_vector(0 downto 0);
      accessReg_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
      accessReg_request_pipe_read_data : in   std_logic_vector(63 downto 0);
      accessReg_response1_pipe_write_req : out  std_logic_vector(0 downto 0);
      accessReg_response1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      accessReg_response1_pipe_write_data : out  std_logic_vector(31 downto 0);
      accessReg_response2_pipe_write_req : out  std_logic_vector(0 downto 0);
      accessReg_response2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      accessReg_response2_pipe_write_data : out  std_logic_vector(31 downto 0);
      accessReg_call_reqs : out  std_logic_vector(0 downto 0);
      accessReg_call_acks : in   std_logic_vector(0 downto 0);
      accessReg_call_data : out  std_logic_vector(58 downto 0);
      accessReg_call_tag  :  out  std_logic_vector(0 downto 0);
      accessReg_return_reqs : out  std_logic_vector(0 downto 0);
      accessReg_return_acks : in   std_logic_vector(0 downto 0);
      accessReg_return_data : in   std_logic_vector(63 downto 0);
      accessReg_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module regAccessDaemon
  signal regAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal regAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal regAccessDaemon_start_req : std_logic;
  signal regAccessDaemon_start_ack : std_logic;
  signal regAccessDaemon_fin_req   : std_logic;
  signal regAccessDaemon_fin_ack : std_logic;
  -- declarations related to module scoreBoard
  -- aggregate signals for read from pipe accessMem_request
  signal accessMem_request_pipe_read_data: std_logic_vector(63 downto 0);
  signal accessMem_request_pipe_read_req: std_logic_vector(0 downto 0);
  signal accessMem_request_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe accessMem_response
  signal accessMem_response_pipe_write_data: std_logic_vector(31 downto 0);
  signal accessMem_response_pipe_write_req: std_logic_vector(0 downto 0);
  signal accessMem_response_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe accessReg_request
  signal accessReg_request_pipe_read_data: std_logic_vector(63 downto 0);
  signal accessReg_request_pipe_read_req: std_logic_vector(0 downto 0);
  signal accessReg_request_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe accessReg_response1
  signal accessReg_response1_pipe_write_data: std_logic_vector(31 downto 0);
  signal accessReg_response1_pipe_write_req: std_logic_vector(0 downto 0);
  signal accessReg_response1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe accessReg_response2
  signal accessReg_response2_pipe_write_data: std_logic_vector(31 downto 0);
  signal accessReg_response2_pipe_write_req: std_logic_vector(0 downto 0);
  signal accessReg_response2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe processor_result
  signal processor_result_pipe_write_data: std_logic_vector(31 downto 0);
  signal processor_result_pipe_write_req: std_logic_vector(0 downto 0);
  signal processor_result_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe start_processor
  signal start_processor_pipe_read_data: std_logic_vector(7 downto 0);
  signal start_processor_pipe_read_req: std_logic_vector(0 downto 0);
  signal start_processor_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module accessMem
  accessMem_read_write_bar <= accessMem_in_args(42 downto 42);
  accessMem_addr <= accessMem_in_args(41 downto 32);
  accessMem_write_data <= accessMem_in_args(31 downto 0);
  accessMem_out_args <= accessMem_read_data ;
  -- call arbiter for module accessMem
  accessMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 43,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessMem_call_reqs,
      call_acks => accessMem_call_acks,
      return_reqs => accessMem_return_reqs,
      return_acks => accessMem_return_acks,
      call_data  => accessMem_call_data,
      call_tag  => accessMem_call_tag,
      return_tag  => accessMem_return_tag,
      call_mtag => accessMem_tag_in,
      return_mtag => accessMem_tag_out,
      return_data =>accessMem_return_data,
      call_mreq => accessMem_start_req,
      call_mack => accessMem_start_ack,
      return_mreq => accessMem_fin_req,
      return_mack => accessMem_fin_ack,
      call_mdata => accessMem_in_args,
      return_mdata => accessMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMem_instance:accessMem-- 
    generic map(tag_length => 4)
    port map(-- 
      read_write_bar => accessMem_read_write_bar,
      addr => accessMem_addr,
      write_data => accessMem_write_data,
      read_data => accessMem_read_data,
      start_req => accessMem_start_req,
      start_ack => accessMem_start_ack,
      fin_req => accessMem_fin_req,
      fin_ack => accessMem_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(9 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(9 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => accessMem_tag_in,
      tag_out => accessMem_tag_out-- 
    ); -- 
  -- module accessReg
  accessReg_valid_1 <= accessReg_in_args(58 downto 58);
  accessReg_addr_1 <= accessReg_in_args(57 downto 50);
  accessReg_valid_2 <= accessReg_in_args(49 downto 49);
  accessReg_addr_2 <= accessReg_in_args(48 downto 41);
  accessReg_valid_w <= accessReg_in_args(40 downto 40);
  accessReg_addr_w <= accessReg_in_args(39 downto 32);
  accessReg_data_to_be_written <= accessReg_in_args(31 downto 0);
  accessReg_out_args <= accessReg_read_data_1 & accessReg_read_data_2 ;
  -- call arbiter for module accessReg
  accessReg_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 59,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessReg_call_reqs,
      call_acks => accessReg_call_acks,
      return_reqs => accessReg_return_reqs,
      return_acks => accessReg_return_acks,
      call_data  => accessReg_call_data,
      call_tag  => accessReg_call_tag,
      return_tag  => accessReg_return_tag,
      call_mtag => accessReg_tag_in,
      return_mtag => accessReg_tag_out,
      return_data =>accessReg_return_data,
      call_mreq => accessReg_start_req,
      call_mack => accessReg_start_ack,
      return_mreq => accessReg_fin_req,
      return_mack => accessReg_fin_ack,
      call_mdata => accessReg_in_args,
      return_mdata => accessReg_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessReg_instance:accessReg-- 
    generic map(tag_length => 3)
    port map(-- 
      valid_1 => accessReg_valid_1,
      addr_1 => accessReg_addr_1,
      valid_2 => accessReg_valid_2,
      addr_2 => accessReg_addr_2,
      valid_w => accessReg_valid_w,
      addr_w => accessReg_addr_w,
      data_to_be_written => accessReg_data_to_be_written,
      read_data_1 => accessReg_read_data_1,
      read_data_2 => accessReg_read_data_2,
      start_req => accessReg_start_req,
      start_ack => accessReg_start_ack,
      fin_req => accessReg_fin_req,
      fin_ack => accessReg_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(5 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(5 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      tag_in => accessReg_tag_in,
      tag_out => accessReg_tag_out-- 
    ); -- 
  -- module iExecStage
  iExecStage_iexec_state <= iExecStage_in_args(169 downto 64);
  iExecStage_iexec_rd1_final <= iExecStage_in_args(63 downto 32);
  iExecStage_iexec_rd2_final <= iExecStage_in_args(31 downto 0);
  iExecStage_out_args <= iExecStage_next_dcache_state ;
  -- call arbiter for module iExecStage
  iExecStage_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 170,
      return_data_width => 139,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => iExecStage_call_reqs,
      call_acks => iExecStage_call_acks,
      return_reqs => iExecStage_return_reqs,
      return_acks => iExecStage_return_acks,
      call_data  => iExecStage_call_data,
      call_tag  => iExecStage_call_tag,
      return_tag  => iExecStage_return_tag,
      call_mtag => iExecStage_tag_in,
      return_mtag => iExecStage_tag_out,
      return_data =>iExecStage_return_data,
      call_mreq => iExecStage_start_req,
      call_mack => iExecStage_start_ack,
      return_mreq => iExecStage_fin_req,
      return_mack => iExecStage_fin_ack,
      call_mdata => iExecStage_in_args,
      return_mdata => iExecStage_out_args,
      clk => clk, 
      reset => reset --
    ); --
  iExecStage_instance:iExecStage-- 
    generic map(tag_length => 2)
    port map(-- 
      iexec_state => iExecStage_iexec_state,
      iexec_rd1_final => iExecStage_iexec_rd1_final,
      iexec_rd2_final => iExecStage_iexec_rd2_final,
      next_dcache_state => iExecStage_next_dcache_state,
      start_req => iExecStage_start_req,
      start_ack => iExecStage_start_ack,
      fin_req => iExecStage_fin_req,
      fin_ack => iExecStage_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => iExecStage_tag_in,
      tag_out => iExecStage_tag_out-- 
    ); -- 
  -- module memAccessDaemon
  memAccessDaemon_instance:memAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => memAccessDaemon_start_req,
      start_ack => memAccessDaemon_start_ack,
      fin_req => memAccessDaemon_fin_req,
      fin_ack => memAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      accessMem_request_pipe_read_req => accessMem_request_pipe_read_req(0 downto 0),
      accessMem_request_pipe_read_ack => accessMem_request_pipe_read_ack(0 downto 0),
      accessMem_request_pipe_read_data => accessMem_request_pipe_read_data(63 downto 0),
      accessMem_response_pipe_write_req => accessMem_response_pipe_write_req(0 downto 0),
      accessMem_response_pipe_write_ack => accessMem_response_pipe_write_ack(0 downto 0),
      accessMem_response_pipe_write_data => accessMem_response_pipe_write_data(31 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(1 downto 1),
      accessMem_call_acks => accessMem_call_acks(1 downto 1),
      accessMem_call_data => accessMem_call_data(85 downto 43),
      accessMem_call_tag => accessMem_call_tag(3 downto 2),
      accessMem_return_reqs => accessMem_return_reqs(1 downto 1),
      accessMem_return_acks => accessMem_return_acks(1 downto 1),
      accessMem_return_data => accessMem_return_data(63 downto 32),
      accessMem_return_tag => accessMem_return_tag(3 downto 2),
      tag_in => memAccessDaemon_tag_in,
      tag_out => memAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  memAccessDaemon_tag_in <= (others => '0');
  memAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => memAccessDaemon_start_req, start_ack => memAccessDaemon_start_ack,  fin_req => memAccessDaemon_fin_req,  fin_ack => memAccessDaemon_fin_ack);
  -- module processor_daemon
  processor_daemon_instance:processor_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => processor_daemon_start_req,
      start_ack => processor_daemon_start_ack,
      fin_req => processor_daemon_fin_req,
      fin_ack => processor_daemon_fin_ack,
      clk => clk,
      reset => reset,
      start_processor_pipe_read_req => start_processor_pipe_read_req(0 downto 0),
      start_processor_pipe_read_ack => start_processor_pipe_read_ack(0 downto 0),
      start_processor_pipe_read_data => start_processor_pipe_read_data(7 downto 0),
      processor_result_pipe_write_req => processor_result_pipe_write_req(0 downto 0),
      processor_result_pipe_write_ack => processor_result_pipe_write_ack(0 downto 0),
      processor_result_pipe_write_data => processor_result_pipe_write_data(31 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(0 downto 0),
      accessMem_call_acks => accessMem_call_acks(0 downto 0),
      accessMem_call_data => accessMem_call_data(42 downto 0),
      accessMem_call_tag => accessMem_call_tag(1 downto 0),
      accessMem_return_reqs => accessMem_return_reqs(0 downto 0),
      accessMem_return_acks => accessMem_return_acks(0 downto 0),
      accessMem_return_data => accessMem_return_data(31 downto 0),
      accessMem_return_tag => accessMem_return_tag(1 downto 0),
      accessReg_call_reqs => accessReg_call_reqs(1 downto 1),
      accessReg_call_acks => accessReg_call_acks(1 downto 1),
      accessReg_call_data => accessReg_call_data(117 downto 59),
      accessReg_call_tag => accessReg_call_tag(1 downto 1),
      accessReg_return_reqs => accessReg_return_reqs(1 downto 1),
      accessReg_return_acks => accessReg_return_acks(1 downto 1),
      accessReg_return_data => accessReg_return_data(127 downto 64),
      accessReg_return_tag => accessReg_return_tag(1 downto 1),
      iExecStage_call_reqs => iExecStage_call_reqs(0 downto 0),
      iExecStage_call_acks => iExecStage_call_acks(0 downto 0),
      iExecStage_call_data => iExecStage_call_data(169 downto 0),
      iExecStage_call_tag => iExecStage_call_tag(0 downto 0),
      iExecStage_return_reqs => iExecStage_return_reqs(0 downto 0),
      iExecStage_return_acks => iExecStage_return_acks(0 downto 0),
      iExecStage_return_data => iExecStage_return_data(138 downto 0),
      iExecStage_return_tag => iExecStage_return_tag(0 downto 0),
      tag_in => processor_daemon_tag_in,
      tag_out => processor_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  processor_daemon_tag_in <= (others => '0');
  processor_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => processor_daemon_start_req, start_ack => processor_daemon_start_ack,  fin_req => processor_daemon_fin_req,  fin_ack => processor_daemon_fin_ack);
  -- module regAccessDaemon
  regAccessDaemon_instance:regAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => regAccessDaemon_start_req,
      start_ack => regAccessDaemon_start_ack,
      fin_req => regAccessDaemon_fin_req,
      fin_ack => regAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      accessReg_request_pipe_read_req => accessReg_request_pipe_read_req(0 downto 0),
      accessReg_request_pipe_read_ack => accessReg_request_pipe_read_ack(0 downto 0),
      accessReg_request_pipe_read_data => accessReg_request_pipe_read_data(63 downto 0),
      accessReg_response1_pipe_write_req => accessReg_response1_pipe_write_req(0 downto 0),
      accessReg_response1_pipe_write_ack => accessReg_response1_pipe_write_ack(0 downto 0),
      accessReg_response1_pipe_write_data => accessReg_response1_pipe_write_data(31 downto 0),
      accessReg_response2_pipe_write_req => accessReg_response2_pipe_write_req(0 downto 0),
      accessReg_response2_pipe_write_ack => accessReg_response2_pipe_write_ack(0 downto 0),
      accessReg_response2_pipe_write_data => accessReg_response2_pipe_write_data(31 downto 0),
      accessReg_call_reqs => accessReg_call_reqs(0 downto 0),
      accessReg_call_acks => accessReg_call_acks(0 downto 0),
      accessReg_call_data => accessReg_call_data(58 downto 0),
      accessReg_call_tag => accessReg_call_tag(0 downto 0),
      accessReg_return_reqs => accessReg_return_reqs(0 downto 0),
      accessReg_return_acks => accessReg_return_acks(0 downto 0),
      accessReg_return_data => accessReg_return_data(63 downto 0),
      accessReg_return_tag => accessReg_return_tag(0 downto 0),
      tag_in => regAccessDaemon_tag_in,
      tag_out => regAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  regAccessDaemon_tag_in <= (others => '0');
  regAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => regAccessDaemon_start_req, start_ack => regAccessDaemon_start_ack,  fin_req => regAccessDaemon_fin_req,  fin_ack => regAccessDaemon_fin_ack);
  accessMem_request_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe accessMem_request",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => accessMem_request_pipe_read_req,
      read_ack => accessMem_request_pipe_read_ack,
      read_data => accessMem_request_pipe_read_data,
      write_req => accessMem_request_pipe_write_req,
      write_ack => accessMem_request_pipe_write_ack,
      write_data => accessMem_request_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  accessMem_response_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe accessMem_response",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => accessMem_response_pipe_read_req,
      read_ack => accessMem_response_pipe_read_ack,
      read_data => accessMem_response_pipe_read_data,
      write_req => accessMem_response_pipe_write_req,
      write_ack => accessMem_response_pipe_write_ack,
      write_data => accessMem_response_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  accessReg_request_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe accessReg_request",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => accessReg_request_pipe_read_req,
      read_ack => accessReg_request_pipe_read_ack,
      read_data => accessReg_request_pipe_read_data,
      write_req => accessReg_request_pipe_write_req,
      write_ack => accessReg_request_pipe_write_ack,
      write_data => accessReg_request_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  accessReg_response1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe accessReg_response1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => accessReg_response1_pipe_read_req,
      read_ack => accessReg_response1_pipe_read_ack,
      read_data => accessReg_response1_pipe_read_data,
      write_req => accessReg_response1_pipe_write_req,
      write_ack => accessReg_response1_pipe_write_ack,
      write_data => accessReg_response1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  accessReg_response2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe accessReg_response2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => accessReg_response2_pipe_read_req,
      read_ack => accessReg_response2_pipe_read_ack,
      read_data => accessReg_response2_pipe_read_data,
      write_req => accessReg_response2_pipe_write_req,
      write_ack => accessReg_response2_pipe_write_ack,
      write_data => accessReg_response2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  processor_result_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe processor_result",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => processor_result_pipe_read_req,
      read_ack => processor_result_pipe_read_ack,
      read_data => processor_result_pipe_read_data,
      write_req => processor_result_pipe_write_req,
      write_ack => processor_result_pipe_write_ack,
      write_data => processor_result_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  start_processor_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe start_processor",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => start_processor_pipe_read_req,
      read_ack => start_processor_pipe_read_ack,
      read_data => start_processor_pipe_read_data,
      write_req => start_processor_pipe_write_req,
      write_ack => start_processor_pipe_write_ack,
      write_data => start_processor_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 10,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 6,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 6,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
